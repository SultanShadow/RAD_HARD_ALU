magic
tech sky130A
magscale 1 2
timestamp 1641133681
<< metal1 >>
rect 198642 700544 198648 700596
rect 198700 700584 198706 700596
rect 283834 700584 283840 700596
rect 198700 700556 283840 700584
rect 198700 700544 198706 700556
rect 283834 700544 283840 700556
rect 283892 700544 283898 700596
rect 206922 700476 206928 700528
rect 206980 700516 206986 700528
rect 348786 700516 348792 700528
rect 206980 700488 348792 700516
rect 206980 700476 206986 700488
rect 348786 700476 348792 700488
rect 348844 700476 348850 700528
rect 249702 700408 249708 700460
rect 249760 700448 249766 700460
rect 413646 700448 413652 700460
rect 249760 700420 413652 700448
rect 249760 700408 249766 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 251818 700340 251824 700392
rect 251876 700380 251882 700392
rect 478506 700380 478512 700392
rect 251876 700352 478512 700380
rect 251876 700340 251882 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 198550 700272 198556 700324
rect 198608 700312 198614 700324
rect 543458 700312 543464 700324
rect 198608 700284 543464 700312
rect 198608 700272 198614 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 198458 683136 198464 683188
rect 198516 683176 198522 683188
rect 580166 683176 580172 683188
rect 198516 683148 580172 683176
rect 198516 683136 198522 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 238662 630640 238668 630692
rect 238720 630680 238726 630692
rect 580166 630680 580172 630692
rect 238720 630652 580172 630680
rect 238720 630640 238726 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 198366 524424 198372 524476
rect 198424 524464 198430 524476
rect 580166 524464 580172 524476
rect 198424 524436 580172 524464
rect 198424 524424 198430 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 234522 470568 234528 470620
rect 234580 470608 234586 470620
rect 580166 470608 580172 470620
rect 234580 470580 580172 470608
rect 234580 470568 234586 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 251910 418140 251916 418192
rect 251968 418180 251974 418192
rect 580166 418180 580172 418192
rect 251968 418152 580172 418180
rect 251968 418140 251974 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 198826 364352 198832 364404
rect 198884 364392 198890 364404
rect 579614 364392 579620 364404
rect 198884 364364 579620 364392
rect 198884 364352 198890 364364
rect 579614 364352 579620 364364
rect 579672 364352 579678 364404
rect 252002 311856 252008 311908
rect 252060 311896 252066 311908
rect 579982 311896 579988 311908
rect 252060 311868 579988 311896
rect 252060 311856 252066 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 198182 258068 198188 258120
rect 198240 258108 198246 258120
rect 580166 258108 580172 258120
rect 198240 258080 580172 258108
rect 198240 258068 198246 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 205818 254736 205824 254788
rect 205876 254776 205882 254788
rect 206922 254776 206928 254788
rect 205876 254748 206928 254776
rect 205876 254736 205882 254748
rect 206922 254736 206928 254748
rect 206980 254736 206986 254788
rect 233510 254736 233516 254788
rect 233568 254776 233574 254788
rect 234522 254776 234528 254788
rect 233568 254748 234528 254776
rect 233568 254736 233574 254748
rect 234522 254736 234528 254748
rect 234580 254736 234586 254788
rect 3418 254668 3424 254720
rect 3476 254708 3482 254720
rect 216766 254708 216772 254720
rect 3476 254680 216772 254708
rect 3476 254668 3482 254680
rect 216766 254668 216772 254680
rect 216824 254668 216830 254720
rect 3602 254600 3608 254652
rect 3660 254640 3666 254652
rect 221918 254640 221924 254652
rect 3660 254612 221924 254640
rect 3660 254600 3666 254612
rect 221918 254600 221924 254612
rect 221976 254600 221982 254652
rect 3878 254532 3884 254584
rect 3936 254572 3942 254584
rect 244458 254572 244464 254584
rect 3936 254544 244464 254572
rect 3936 254532 3942 254544
rect 244458 254532 244464 254544
rect 244516 254532 244522 254584
rect 2682 253920 2688 253972
rect 2740 253960 2746 253972
rect 200022 253960 200028 253972
rect 2740 253932 200028 253960
rect 2740 253920 2746 253932
rect 200022 253920 200028 253932
rect 200080 253920 200086 253972
rect 227714 253920 227720 253972
rect 227772 253960 227778 253972
rect 250438 253960 250444 253972
rect 227772 253932 250444 253960
rect 227772 253920 227778 253932
rect 250438 253920 250444 253932
rect 250496 253920 250502 253972
rect 89622 241408 89628 241460
rect 89680 241448 89686 241460
rect 197906 241448 197912 241460
rect 89680 241420 197912 241448
rect 89680 241408 89686 241420
rect 197906 241408 197912 241420
rect 197964 241408 197970 241460
rect 3694 223524 3700 223576
rect 3752 223564 3758 223576
rect 197354 223564 197360 223576
rect 3752 223536 197360 223564
rect 3752 223524 3758 223536
rect 197354 223524 197360 223536
rect 197412 223524 197418 223576
rect 3142 202036 3148 202088
rect 3200 202076 3206 202088
rect 251174 202076 251180 202088
rect 3200 202048 251180 202076
rect 3200 202036 3206 202048
rect 251174 202036 251180 202048
rect 251232 202036 251238 202088
rect 3970 198636 3976 198688
rect 4028 198676 4034 198688
rect 210970 198676 210976 198688
rect 4028 198648 210976 198676
rect 4028 198636 4034 198648
rect 210970 198636 210976 198648
rect 211028 198636 211034 198688
rect 216122 198636 216128 198688
rect 216180 198676 216186 198688
rect 580258 198676 580264 198688
rect 216180 198648 580264 198676
rect 216180 198636 216186 198648
rect 580258 198636 580264 198648
rect 580316 198636 580322 198688
rect 3786 198568 3792 198620
rect 3844 198608 3850 198620
rect 238662 198608 238668 198620
rect 3844 198580 238668 198608
rect 3844 198568 3850 198580
rect 238662 198568 238668 198580
rect 238720 198568 238726 198620
rect 249610 198568 249616 198620
rect 249668 198608 249674 198620
rect 580350 198608 580356 198620
rect 249668 198580 580356 198608
rect 249668 198568 249674 198580
rect 580350 198568 580356 198580
rect 580408 198568 580414 198620
rect 3510 198500 3516 198552
rect 3568 198540 3574 198552
rect 232866 198540 232872 198552
rect 3568 198512 232872 198540
rect 3568 198500 3574 198512
rect 232866 198500 232872 198512
rect 232924 198500 232930 198552
rect 3878 198432 3884 198484
rect 3936 198472 3942 198484
rect 205174 198472 205180 198484
rect 3936 198444 205180 198472
rect 3936 198432 3942 198444
rect 205174 198432 205180 198444
rect 205232 198432 205238 198484
rect 154482 198364 154488 198416
rect 154540 198404 154546 198416
rect 221918 198404 221924 198416
rect 154540 198376 221924 198404
rect 154540 198364 154546 198376
rect 221918 198364 221924 198376
rect 221976 198364 221982 198416
rect 227714 197888 227720 197940
rect 227772 197928 227778 197940
rect 229002 197928 229008 197940
rect 227772 197900 229008 197928
rect 227772 197888 227778 197900
rect 229002 197888 229008 197900
rect 229060 197888 229066 197940
rect 198274 179324 198280 179376
rect 198332 179364 198338 179376
rect 580166 179364 580172 179376
rect 198332 179336 580172 179364
rect 198332 179324 198338 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 250438 139340 250444 139392
rect 250496 139380 250502 139392
rect 580166 139380 580172 139392
rect 250496 139352 580172 139380
rect 250496 139340 250502 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 229002 100648 229008 100700
rect 229060 100688 229066 100700
rect 580166 100688 580172 100700
rect 229060 100660 580172 100688
rect 229060 100648 229066 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 251818 46860 251824 46912
rect 251876 46900 251882 46912
rect 580166 46900 580172 46912
rect 251876 46872 580172 46900
rect 251876 46860 251882 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 244182 3408 244188 3460
rect 244240 3448 244246 3460
rect 579798 3448 579804 3460
rect 244240 3420 579804 3448
rect 244240 3408 244246 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
<< via1 >>
rect 198648 700544 198700 700596
rect 283840 700544 283892 700596
rect 206928 700476 206980 700528
rect 348792 700476 348844 700528
rect 249708 700408 249760 700460
rect 413652 700408 413704 700460
rect 251824 700340 251876 700392
rect 478512 700340 478564 700392
rect 198556 700272 198608 700324
rect 543464 700272 543516 700324
rect 198464 683136 198516 683188
rect 580172 683136 580224 683188
rect 238668 630640 238720 630692
rect 580172 630640 580224 630692
rect 198372 524424 198424 524476
rect 580172 524424 580224 524476
rect 234528 470568 234580 470620
rect 580172 470568 580224 470620
rect 251916 418140 251968 418192
rect 580172 418140 580224 418192
rect 198832 364352 198884 364404
rect 579620 364352 579672 364404
rect 252008 311856 252060 311908
rect 579988 311856 580040 311908
rect 198188 258068 198240 258120
rect 580172 258068 580224 258120
rect 205824 254736 205876 254788
rect 206928 254736 206980 254788
rect 233516 254736 233568 254788
rect 234528 254736 234580 254788
rect 3424 254668 3476 254720
rect 216772 254668 216824 254720
rect 3608 254600 3660 254652
rect 221924 254600 221976 254652
rect 3884 254532 3936 254584
rect 244464 254532 244516 254584
rect 2688 253920 2740 253972
rect 200028 253920 200080 253972
rect 227720 253920 227772 253972
rect 250444 253920 250496 253972
rect 89628 241408 89680 241460
rect 197912 241408 197964 241460
rect 3700 223524 3752 223576
rect 197360 223524 197412 223576
rect 3148 202036 3200 202088
rect 251180 202036 251232 202088
rect 3976 198636 4028 198688
rect 210976 198636 211028 198688
rect 216128 198636 216180 198688
rect 580264 198636 580316 198688
rect 3792 198568 3844 198620
rect 238668 198568 238720 198620
rect 249616 198568 249668 198620
rect 580356 198568 580408 198620
rect 3516 198500 3568 198552
rect 232872 198500 232924 198552
rect 3884 198432 3936 198484
rect 205180 198432 205232 198484
rect 154488 198364 154540 198416
rect 221924 198364 221976 198416
rect 227720 197888 227772 197940
rect 229008 197888 229060 197940
rect 198280 179324 198332 179376
rect 580172 179324 580224 179376
rect 250444 139340 250496 139392
rect 580172 139340 580224 139392
rect 229008 100648 229060 100700
rect 580172 100648 580224 100700
rect 251824 46860 251876 46912
rect 580172 46860 580224 46912
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 244188 3408 244240 3460
rect 579804 3408 579856 3460
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 89364 703582 89668 703610
rect 24320 699825 24348 703520
rect 89180 703474 89208 703520
rect 89364 703474 89392 703582
rect 89180 703446 89392 703474
rect 24306 699816 24362 699825
rect 24306 699751 24362 699760
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 254726 3464 671191
rect 3606 619168 3662 619177
rect 3606 619103 3662 619112
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3424 254720 3476 254726
rect 3424 254662 3476 254668
rect 2688 253972 2740 253978
rect 2688 253914 2740 253920
rect 2700 3534 2728 253914
rect 3148 202088 3200 202094
rect 3148 202030 3200 202036
rect 3160 201929 3188 202030
rect 3146 201920 3202 201929
rect 3146 201855 3202 201864
rect 3528 198558 3556 566879
rect 3620 254658 3648 619103
rect 3698 514856 3754 514865
rect 3698 514791 3754 514800
rect 3608 254652 3660 254658
rect 3608 254594 3660 254600
rect 3712 223582 3740 514791
rect 3790 462632 3846 462641
rect 3790 462567 3846 462576
rect 3700 223576 3752 223582
rect 3700 223518 3752 223524
rect 3804 198626 3832 462567
rect 3882 410544 3938 410553
rect 3882 410479 3938 410488
rect 3896 254590 3924 410479
rect 3974 306232 4030 306241
rect 3974 306167 4030 306176
rect 3884 254584 3936 254590
rect 3884 254526 3936 254532
rect 3988 209774 4016 306167
rect 4066 254144 4122 254153
rect 4066 254079 4122 254088
rect 3896 209746 4016 209774
rect 3792 198620 3844 198626
rect 3792 198562 3844 198568
rect 3516 198552 3568 198558
rect 3516 198494 3568 198500
rect 3896 198490 3924 209746
rect 4080 200114 4108 254079
rect 89640 241466 89668 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 154316 703582 154528 703610
rect 154132 703474 154160 703520
rect 154316 703474 154344 703582
rect 154132 703446 154344 703474
rect 89628 241460 89680 241466
rect 89628 241402 89680 241408
rect 3988 200086 4108 200114
rect 3988 198694 4016 200086
rect 3976 198688 4028 198694
rect 3976 198630 4028 198636
rect 3884 198484 3936 198490
rect 3884 198426 3936 198432
rect 154500 198422 154528 703582
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 198648 700596 198700 700602
rect 198648 700538 198700 700544
rect 198556 700324 198608 700330
rect 198556 700266 198608 700272
rect 198464 683188 198516 683194
rect 198464 683130 198516 683136
rect 198372 524476 198424 524482
rect 198372 524418 198424 524424
rect 198188 258120 198240 258126
rect 198188 258062 198240 258068
rect 197912 241460 197964 241466
rect 197912 241402 197964 241408
rect 197924 240961 197952 241402
rect 197910 240952 197966 240961
rect 197910 240887 197966 240896
rect 197360 223576 197412 223582
rect 197360 223518 197412 223524
rect 197372 223281 197400 223518
rect 197358 223272 197414 223281
rect 197358 223207 197414 223216
rect 198200 205601 198228 258062
rect 198278 246392 198334 246401
rect 198278 246327 198334 246336
rect 198186 205592 198242 205601
rect 198186 205527 198242 205536
rect 154488 198416 154540 198422
rect 154488 198358 154540 198364
rect 198292 179382 198320 246327
rect 198384 234841 198412 524418
rect 198370 234832 198426 234841
rect 198370 234767 198426 234776
rect 198476 217161 198504 683130
rect 198568 229401 198596 700266
rect 198554 229392 198610 229401
rect 198554 229327 198610 229336
rect 198462 217152 198518 217161
rect 198462 217087 198518 217096
rect 198660 211721 198688 700538
rect 206928 700528 206980 700534
rect 206928 700470 206980 700476
rect 198832 364404 198884 364410
rect 198832 364346 198884 364352
rect 198646 211712 198702 211721
rect 198646 211647 198702 211656
rect 198844 209774 198872 364346
rect 206940 254794 206968 700470
rect 218992 699825 219020 703520
rect 283852 700602 283880 703520
rect 283840 700596 283892 700602
rect 283840 700538 283892 700544
rect 348804 700534 348832 703520
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 413664 700466 413692 703520
rect 249708 700460 249760 700466
rect 249708 700402 249760 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 218978 699816 219034 699825
rect 218978 699751 219034 699760
rect 238668 630692 238720 630698
rect 238668 630634 238720 630640
rect 234528 470620 234580 470626
rect 234528 470562 234580 470568
rect 234540 254794 234568 470562
rect 205824 254788 205876 254794
rect 205824 254730 205876 254736
rect 206928 254788 206980 254794
rect 206928 254730 206980 254736
rect 233516 254788 233568 254794
rect 233516 254730 233568 254736
rect 234528 254788 234580 254794
rect 234528 254730 234580 254736
rect 200028 253972 200080 253978
rect 200028 253914 200080 253920
rect 200040 252212 200068 253914
rect 205836 252212 205864 254730
rect 216772 254720 216824 254726
rect 216772 254662 216824 254668
rect 216784 252212 216812 254662
rect 221924 254652 221976 254658
rect 221924 254594 221976 254600
rect 221936 252212 221964 254594
rect 227720 253972 227772 253978
rect 227720 253914 227772 253920
rect 227732 252212 227760 253914
rect 233528 252212 233556 254730
rect 238680 252212 238708 630634
rect 244464 254584 244516 254590
rect 244464 254526 244516 254532
rect 244476 252212 244504 254526
rect 249720 252226 249748 700402
rect 478524 700398 478552 703520
rect 251824 700392 251876 700398
rect 251824 700334 251876 700340
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 250444 253972 250496 253978
rect 250444 253914 250496 253920
rect 249642 252198 249748 252226
rect 210698 251696 210754 251705
rect 210754 251654 211002 251682
rect 210698 251631 210754 251640
rect 198844 209746 199608 209774
rect 199580 200682 199608 209746
rect 199580 200654 200054 200682
rect 205192 198490 205220 200124
rect 210988 198694 211016 200124
rect 216140 198694 216168 200124
rect 210976 198688 211028 198694
rect 210976 198630 211028 198636
rect 216128 198688 216180 198694
rect 216128 198630 216180 198636
rect 205180 198484 205232 198490
rect 205180 198426 205232 198432
rect 221936 198422 221964 200124
rect 221924 198416 221976 198422
rect 221924 198358 221976 198364
rect 227732 197946 227760 200124
rect 232884 198558 232912 200124
rect 238680 198626 238708 200124
rect 243846 200110 244228 200138
rect 238668 198620 238720 198626
rect 238668 198562 238720 198568
rect 232872 198552 232924 198558
rect 232872 198494 232924 198500
rect 227720 197940 227772 197946
rect 227720 197882 227772 197888
rect 229008 197940 229060 197946
rect 229008 197882 229060 197888
rect 198280 179376 198332 179382
rect 198280 179318 198332 179324
rect 229020 100706 229048 197882
rect 229008 100700 229060 100706
rect 229008 100642 229060 100648
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 1688 480 1716 3470
rect 244200 3466 244228 200110
rect 249628 198626 249656 200124
rect 249616 198620 249668 198626
rect 249616 198562 249668 198568
rect 250456 139398 250484 253914
rect 251178 240408 251234 240417
rect 251178 240343 251234 240352
rect 251192 202094 251220 240343
rect 251836 228857 251864 700334
rect 543476 700330 543504 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 251916 418192 251968 418198
rect 251916 418134 251968 418140
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 251822 228848 251878 228857
rect 251822 228783 251878 228792
rect 251822 222320 251878 222329
rect 251822 222255 251878 222264
rect 251180 202088 251232 202094
rect 251180 202030 251232 202036
rect 250444 139392 250496 139398
rect 250444 139334 250496 139340
rect 251836 46918 251864 222255
rect 251928 211177 251956 418134
rect 579618 365120 579674 365129
rect 579618 365055 579674 365064
rect 579632 364410 579660 365055
rect 579620 364404 579672 364410
rect 579620 364346 579672 364352
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 252008 311908 252060 311914
rect 252008 311850 252060 311856
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 252020 235385 252048 311850
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 252006 235376 252062 235385
rect 252006 235311 252062 235320
rect 251914 211168 251970 211177
rect 251914 211103 251970 211112
rect 580276 198694 580304 577623
rect 580354 219056 580410 219065
rect 580354 218991 580410 219000
rect 580264 198688 580316 198694
rect 580264 198630 580316 198636
rect 580368 198626 580396 218991
rect 580356 198620 580408 198626
rect 580356 198562 580408 198568
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 251824 46912 251876 46918
rect 251824 46854 251876 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 244188 3460 244240 3466
rect 244188 3402 244240 3408
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 24306 699760 24362 699816
rect 3422 671200 3478 671256
rect 3606 619112 3662 619168
rect 3514 566888 3570 566944
rect 3146 201864 3202 201920
rect 3698 514800 3754 514856
rect 3790 462576 3846 462632
rect 3882 410488 3938 410544
rect 3974 306176 4030 306232
rect 4066 254088 4122 254144
rect 197910 240896 197966 240952
rect 197358 223216 197414 223272
rect 198278 246336 198334 246392
rect 198186 205536 198242 205592
rect 198370 234776 198426 234832
rect 198554 229336 198610 229392
rect 198462 217096 198518 217152
rect 198646 211656 198702 211712
rect 218978 699760 219034 699816
rect 210698 251640 210754 251696
rect 251178 240352 251234 240408
rect 580170 683848 580226 683904
rect 580170 630808 580226 630864
rect 580262 577632 580318 577688
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 471416 580226 471472
rect 580170 418240 580226 418296
rect 251822 228792 251878 228848
rect 251822 222264 251878 222320
rect 579618 365064 579674 365120
rect 579986 312024 580042 312080
rect 580170 258848 580226 258904
rect 252006 235320 252062 235376
rect 251914 211112 251970 211168
rect 580354 219000 580410 219056
rect 580170 179152 580226 179208
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 99456 580226 99512
rect 580170 46280 580226 46336
<< metal3 >>
rect 24301 699818 24367 699821
rect 24710 699818 24716 699820
rect 24301 699816 24716 699818
rect 24301 699760 24306 699816
rect 24362 699760 24716 699816
rect 24301 699758 24716 699760
rect 24301 699755 24367 699758
rect 24710 699756 24716 699758
rect 24780 699756 24786 699820
rect 218973 699818 219039 699821
rect 219198 699818 219204 699820
rect 218973 699816 219204 699818
rect 218973 699760 218978 699816
rect 219034 699760 219204 699816
rect 218973 699758 219204 699760
rect 218973 699755 219039 699758
rect 219198 699756 219204 699758
rect 219268 699756 219274 699820
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3601 619170 3667 619173
rect -960 619168 3667 619170
rect -960 619112 3606 619168
rect 3662 619112 3667 619168
rect -960 619110 3667 619112
rect -960 619020 480 619110
rect 3601 619107 3667 619110
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3693 514858 3759 514861
rect -960 514856 3759 514858
rect -960 514800 3698 514856
rect 3754 514800 3759 514856
rect -960 514798 3759 514800
rect -960 514708 480 514798
rect 3693 514795 3759 514798
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3785 462634 3851 462637
rect -960 462632 3851 462634
rect -960 462576 3790 462632
rect 3846 462576 3851 462632
rect -960 462574 3851 462576
rect -960 462484 480 462574
rect 3785 462571 3851 462574
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3877 410546 3943 410549
rect -960 410544 3943 410546
rect -960 410488 3882 410544
rect 3938 410488 3943 410544
rect -960 410486 3943 410488
rect -960 410396 480 410486
rect 3877 410483 3943 410486
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 579613 365122 579679 365125
rect 583520 365122 584960 365212
rect 579613 365120 584960 365122
rect 579613 365064 579618 365120
rect 579674 365064 584960 365120
rect 579613 365062 584960 365064
rect 579613 365059 579679 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3366 358458 3372 358460
rect -960 358398 3372 358458
rect -960 358308 480 358398
rect 3366 358396 3372 358398
rect 3436 358396 3442 358460
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3969 306234 4035 306237
rect -960 306232 4035 306234
rect -960 306176 3974 306232
rect 4030 306176 4035 306232
rect -960 306174 4035 306176
rect -960 306084 480 306174
rect 3969 306171 4035 306174
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 4061 254146 4127 254149
rect -960 254144 4127 254146
rect -960 254088 4066 254144
rect 4122 254088 4127 254144
rect -960 254086 4127 254088
rect -960 253996 480 254086
rect 4061 254083 4127 254086
rect 210550 251636 210556 251700
rect 210620 251698 210626 251700
rect 210693 251698 210759 251701
rect 210620 251696 210759 251698
rect 210620 251640 210698 251696
rect 210754 251640 210759 251696
rect 210620 251638 210759 251640
rect 210620 251636 210626 251638
rect 210693 251635 210759 251638
rect 249558 246876 249564 246940
rect 249628 246876 249634 246940
rect 198273 246394 198339 246397
rect 198273 246392 200100 246394
rect 198273 246336 198278 246392
rect 198334 246336 200100 246392
rect 249566 246364 249626 246876
rect 198273 246334 200100 246336
rect 198273 246331 198339 246334
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 197905 240954 197971 240957
rect 197905 240952 200100 240954
rect 197905 240896 197910 240952
rect 197966 240896 200100 240952
rect 197905 240894 200100 240896
rect 197905 240891 197971 240894
rect 251173 240410 251239 240413
rect 249934 240408 251239 240410
rect 249934 240352 251178 240408
rect 251234 240352 251239 240408
rect 249934 240350 251239 240352
rect 249934 240244 249994 240350
rect 251173 240347 251239 240350
rect 252001 235378 252067 235381
rect 249934 235376 252067 235378
rect 249934 235320 252006 235376
rect 252062 235320 252067 235376
rect 249934 235318 252067 235320
rect 198365 234834 198431 234837
rect 198365 234832 200100 234834
rect 198365 234776 198370 234832
rect 198426 234776 200100 234832
rect 249934 234804 249994 235318
rect 252001 235315 252067 235318
rect 198365 234774 200100 234776
rect 198365 234771 198431 234774
rect 583520 232236 584960 232476
rect 198549 229394 198615 229397
rect 198549 229392 200100 229394
rect 198549 229336 198554 229392
rect 198610 229336 200100 229392
rect 198549 229334 200100 229336
rect 198549 229331 198615 229334
rect 251817 228850 251883 228853
rect 249934 228848 251883 228850
rect 249934 228792 251822 228848
rect 251878 228792 251883 228848
rect 249934 228790 251883 228792
rect 249934 228684 249994 228790
rect 251817 228787 251883 228790
rect -960 227884 480 228124
rect 197353 223274 197419 223277
rect 197353 223272 200100 223274
rect 197353 223216 197358 223272
rect 197414 223216 200100 223272
rect 197353 223214 200100 223216
rect 197353 223211 197419 223214
rect 250118 222322 250178 222564
rect 251817 222322 251883 222325
rect 250118 222320 251883 222322
rect 250118 222264 251822 222320
rect 251878 222264 251883 222320
rect 250118 222262 251883 222264
rect 251817 222259 251883 222262
rect 580349 219058 580415 219061
rect 583520 219058 584960 219148
rect 580349 219056 584960 219058
rect 580349 219000 580354 219056
rect 580410 219000 584960 219056
rect 580349 218998 584960 219000
rect 580349 218995 580415 218998
rect 583520 218908 584960 218998
rect 249558 217636 249564 217700
rect 249628 217636 249634 217700
rect 198457 217154 198523 217157
rect 198457 217152 200100 217154
rect 198457 217096 198462 217152
rect 198518 217096 200100 217152
rect 249566 217124 249626 217636
rect 198457 217094 200100 217096
rect 198457 217091 198523 217094
rect -960 214828 480 215068
rect 198641 211714 198707 211717
rect 198641 211712 200100 211714
rect 198641 211656 198646 211712
rect 198702 211656 200100 211712
rect 198641 211654 200100 211656
rect 198641 211651 198707 211654
rect 251909 211170 251975 211173
rect 249934 211168 251975 211170
rect 249934 211112 251914 211168
rect 251970 211112 251975 211168
rect 249934 211110 251975 211112
rect 249934 211004 249994 211110
rect 251909 211107 251975 211110
rect 198181 205594 198247 205597
rect 198181 205592 200100 205594
rect 198181 205536 198186 205592
rect 198242 205536 200100 205592
rect 583520 205580 584960 205820
rect 198181 205534 200100 205536
rect 198181 205531 198247 205534
rect 249566 205052 249626 205564
rect 249558 204988 249564 205052
rect 249628 204988 249634 205052
rect -960 201922 480 202012
rect 3141 201922 3207 201925
rect -960 201920 3207 201922
rect -960 201864 3146 201920
rect 3202 201864 3207 201920
rect -960 201862 3207 201864
rect -960 201772 480 201862
rect 3141 201859 3207 201862
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect 583520 6626 584960 6716
rect -960 6340 480 6580
rect 583342 6566 584960 6626
rect 583342 6490 583402 6566
rect 583520 6490 584960 6566
rect 583342 6476 584960 6490
rect 583342 6430 583586 6476
rect 210550 5612 210556 5676
rect 210620 5674 210626 5676
rect 583526 5674 583586 6430
rect 210620 5614 583586 5674
rect 210620 5612 210626 5614
<< via3 >>
rect 24716 699756 24780 699820
rect 219204 699756 219268 699820
rect 3372 358396 3436 358460
rect 210556 251636 210620 251700
rect 249564 246876 249628 246940
rect 249564 217636 249628 217700
rect 249564 204988 249628 205052
rect 210556 5612 210620 5676
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 643614 -8106 711002
rect -8726 643378 -8694 643614
rect -8458 643378 -8374 643614
rect -8138 643378 -8106 643614
rect -8726 643294 -8106 643378
rect -8726 643058 -8694 643294
rect -8458 643058 -8374 643294
rect -8138 643058 -8106 643294
rect -8726 583614 -8106 643058
rect -8726 583378 -8694 583614
rect -8458 583378 -8374 583614
rect -8138 583378 -8106 583614
rect -8726 583294 -8106 583378
rect -8726 583058 -8694 583294
rect -8458 583058 -8374 583294
rect -8138 583058 -8106 583294
rect -8726 523614 -8106 583058
rect -8726 523378 -8694 523614
rect -8458 523378 -8374 523614
rect -8138 523378 -8106 523614
rect -8726 523294 -8106 523378
rect -8726 523058 -8694 523294
rect -8458 523058 -8374 523294
rect -8138 523058 -8106 523294
rect -8726 463614 -8106 523058
rect -8726 463378 -8694 463614
rect -8458 463378 -8374 463614
rect -8138 463378 -8106 463614
rect -8726 463294 -8106 463378
rect -8726 463058 -8694 463294
rect -8458 463058 -8374 463294
rect -8138 463058 -8106 463294
rect -8726 403614 -8106 463058
rect -8726 403378 -8694 403614
rect -8458 403378 -8374 403614
rect -8138 403378 -8106 403614
rect -8726 403294 -8106 403378
rect -8726 403058 -8694 403294
rect -8458 403058 -8374 403294
rect -8138 403058 -8106 403294
rect -8726 343614 -8106 403058
rect -8726 343378 -8694 343614
rect -8458 343378 -8374 343614
rect -8138 343378 -8106 343614
rect -8726 343294 -8106 343378
rect -8726 343058 -8694 343294
rect -8458 343058 -8374 343294
rect -8138 343058 -8106 343294
rect -8726 283614 -8106 343058
rect -8726 283378 -8694 283614
rect -8458 283378 -8374 283614
rect -8138 283378 -8106 283614
rect -8726 283294 -8106 283378
rect -8726 283058 -8694 283294
rect -8458 283058 -8374 283294
rect -8138 283058 -8106 283294
rect -8726 223614 -8106 283058
rect -8726 223378 -8694 223614
rect -8458 223378 -8374 223614
rect -8138 223378 -8106 223614
rect -8726 223294 -8106 223378
rect -8726 223058 -8694 223294
rect -8458 223058 -8374 223294
rect -8138 223058 -8106 223294
rect -8726 163614 -8106 223058
rect -8726 163378 -8694 163614
rect -8458 163378 -8374 163614
rect -8138 163378 -8106 163614
rect -8726 163294 -8106 163378
rect -8726 163058 -8694 163294
rect -8458 163058 -8374 163294
rect -8138 163058 -8106 163294
rect -8726 103614 -8106 163058
rect -8726 103378 -8694 103614
rect -8458 103378 -8374 103614
rect -8138 103378 -8106 103614
rect -8726 103294 -8106 103378
rect -8726 103058 -8694 103294
rect -8458 103058 -8374 103294
rect -8138 103058 -8106 103294
rect -8726 43614 -8106 103058
rect -8726 43378 -8694 43614
rect -8458 43378 -8374 43614
rect -8138 43378 -8106 43614
rect -8726 43294 -8106 43378
rect -8726 43058 -8694 43294
rect -8458 43058 -8374 43294
rect -8138 43058 -8106 43294
rect -8726 -7066 -8106 43058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673614 -7146 710042
rect 11954 710598 12574 711590
rect 11954 710362 11986 710598
rect 12222 710362 12306 710598
rect 12542 710362 12574 710598
rect 11954 710278 12574 710362
rect 11954 710042 11986 710278
rect 12222 710042 12306 710278
rect 12542 710042 12574 710278
rect -7766 673378 -7734 673614
rect -7498 673378 -7414 673614
rect -7178 673378 -7146 673614
rect -7766 673294 -7146 673378
rect -7766 673058 -7734 673294
rect -7498 673058 -7414 673294
rect -7178 673058 -7146 673294
rect -7766 613614 -7146 673058
rect -7766 613378 -7734 613614
rect -7498 613378 -7414 613614
rect -7178 613378 -7146 613614
rect -7766 613294 -7146 613378
rect -7766 613058 -7734 613294
rect -7498 613058 -7414 613294
rect -7178 613058 -7146 613294
rect -7766 553614 -7146 613058
rect -7766 553378 -7734 553614
rect -7498 553378 -7414 553614
rect -7178 553378 -7146 553614
rect -7766 553294 -7146 553378
rect -7766 553058 -7734 553294
rect -7498 553058 -7414 553294
rect -7178 553058 -7146 553294
rect -7766 493614 -7146 553058
rect -7766 493378 -7734 493614
rect -7498 493378 -7414 493614
rect -7178 493378 -7146 493614
rect -7766 493294 -7146 493378
rect -7766 493058 -7734 493294
rect -7498 493058 -7414 493294
rect -7178 493058 -7146 493294
rect -7766 433614 -7146 493058
rect -7766 433378 -7734 433614
rect -7498 433378 -7414 433614
rect -7178 433378 -7146 433614
rect -7766 433294 -7146 433378
rect -7766 433058 -7734 433294
rect -7498 433058 -7414 433294
rect -7178 433058 -7146 433294
rect -7766 373614 -7146 433058
rect -7766 373378 -7734 373614
rect -7498 373378 -7414 373614
rect -7178 373378 -7146 373614
rect -7766 373294 -7146 373378
rect -7766 373058 -7734 373294
rect -7498 373058 -7414 373294
rect -7178 373058 -7146 373294
rect -7766 313614 -7146 373058
rect -7766 313378 -7734 313614
rect -7498 313378 -7414 313614
rect -7178 313378 -7146 313614
rect -7766 313294 -7146 313378
rect -7766 313058 -7734 313294
rect -7498 313058 -7414 313294
rect -7178 313058 -7146 313294
rect -7766 253614 -7146 313058
rect -7766 253378 -7734 253614
rect -7498 253378 -7414 253614
rect -7178 253378 -7146 253614
rect -7766 253294 -7146 253378
rect -7766 253058 -7734 253294
rect -7498 253058 -7414 253294
rect -7178 253058 -7146 253294
rect -7766 193614 -7146 253058
rect -7766 193378 -7734 193614
rect -7498 193378 -7414 193614
rect -7178 193378 -7146 193614
rect -7766 193294 -7146 193378
rect -7766 193058 -7734 193294
rect -7498 193058 -7414 193294
rect -7178 193058 -7146 193294
rect -7766 133614 -7146 193058
rect -7766 133378 -7734 133614
rect -7498 133378 -7414 133614
rect -7178 133378 -7146 133614
rect -7766 133294 -7146 133378
rect -7766 133058 -7734 133294
rect -7498 133058 -7414 133294
rect -7178 133058 -7146 133294
rect -7766 73614 -7146 133058
rect -7766 73378 -7734 73614
rect -7498 73378 -7414 73614
rect -7178 73378 -7146 73614
rect -7766 73294 -7146 73378
rect -7766 73058 -7734 73294
rect -7498 73058 -7414 73294
rect -7178 73058 -7146 73294
rect -7766 13614 -7146 73058
rect -7766 13378 -7734 13614
rect -7498 13378 -7414 13614
rect -7178 13378 -7146 13614
rect -7766 13294 -7146 13378
rect -7766 13058 -7734 13294
rect -7498 13058 -7414 13294
rect -7178 13058 -7146 13294
rect -7766 -6106 -7146 13058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 699894 -6186 709082
rect -6806 699658 -6774 699894
rect -6538 699658 -6454 699894
rect -6218 699658 -6186 699894
rect -6806 699574 -6186 699658
rect -6806 699338 -6774 699574
rect -6538 699338 -6454 699574
rect -6218 699338 -6186 699574
rect -6806 639894 -6186 699338
rect -6806 639658 -6774 639894
rect -6538 639658 -6454 639894
rect -6218 639658 -6186 639894
rect -6806 639574 -6186 639658
rect -6806 639338 -6774 639574
rect -6538 639338 -6454 639574
rect -6218 639338 -6186 639574
rect -6806 579894 -6186 639338
rect -6806 579658 -6774 579894
rect -6538 579658 -6454 579894
rect -6218 579658 -6186 579894
rect -6806 579574 -6186 579658
rect -6806 579338 -6774 579574
rect -6538 579338 -6454 579574
rect -6218 579338 -6186 579574
rect -6806 519894 -6186 579338
rect -6806 519658 -6774 519894
rect -6538 519658 -6454 519894
rect -6218 519658 -6186 519894
rect -6806 519574 -6186 519658
rect -6806 519338 -6774 519574
rect -6538 519338 -6454 519574
rect -6218 519338 -6186 519574
rect -6806 459894 -6186 519338
rect -6806 459658 -6774 459894
rect -6538 459658 -6454 459894
rect -6218 459658 -6186 459894
rect -6806 459574 -6186 459658
rect -6806 459338 -6774 459574
rect -6538 459338 -6454 459574
rect -6218 459338 -6186 459574
rect -6806 399894 -6186 459338
rect -6806 399658 -6774 399894
rect -6538 399658 -6454 399894
rect -6218 399658 -6186 399894
rect -6806 399574 -6186 399658
rect -6806 399338 -6774 399574
rect -6538 399338 -6454 399574
rect -6218 399338 -6186 399574
rect -6806 339894 -6186 399338
rect -6806 339658 -6774 339894
rect -6538 339658 -6454 339894
rect -6218 339658 -6186 339894
rect -6806 339574 -6186 339658
rect -6806 339338 -6774 339574
rect -6538 339338 -6454 339574
rect -6218 339338 -6186 339574
rect -6806 279894 -6186 339338
rect -6806 279658 -6774 279894
rect -6538 279658 -6454 279894
rect -6218 279658 -6186 279894
rect -6806 279574 -6186 279658
rect -6806 279338 -6774 279574
rect -6538 279338 -6454 279574
rect -6218 279338 -6186 279574
rect -6806 219894 -6186 279338
rect -6806 219658 -6774 219894
rect -6538 219658 -6454 219894
rect -6218 219658 -6186 219894
rect -6806 219574 -6186 219658
rect -6806 219338 -6774 219574
rect -6538 219338 -6454 219574
rect -6218 219338 -6186 219574
rect -6806 159894 -6186 219338
rect -6806 159658 -6774 159894
rect -6538 159658 -6454 159894
rect -6218 159658 -6186 159894
rect -6806 159574 -6186 159658
rect -6806 159338 -6774 159574
rect -6538 159338 -6454 159574
rect -6218 159338 -6186 159574
rect -6806 99894 -6186 159338
rect -6806 99658 -6774 99894
rect -6538 99658 -6454 99894
rect -6218 99658 -6186 99894
rect -6806 99574 -6186 99658
rect -6806 99338 -6774 99574
rect -6538 99338 -6454 99574
rect -6218 99338 -6186 99574
rect -6806 39894 -6186 99338
rect -6806 39658 -6774 39894
rect -6538 39658 -6454 39894
rect -6218 39658 -6186 39894
rect -6806 39574 -6186 39658
rect -6806 39338 -6774 39574
rect -6538 39338 -6454 39574
rect -6218 39338 -6186 39574
rect -6806 -5146 -6186 39338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669894 -5226 708122
rect 8234 708678 8854 709670
rect 8234 708442 8266 708678
rect 8502 708442 8586 708678
rect 8822 708442 8854 708678
rect 8234 708358 8854 708442
rect 8234 708122 8266 708358
rect 8502 708122 8586 708358
rect 8822 708122 8854 708358
rect -5846 669658 -5814 669894
rect -5578 669658 -5494 669894
rect -5258 669658 -5226 669894
rect -5846 669574 -5226 669658
rect -5846 669338 -5814 669574
rect -5578 669338 -5494 669574
rect -5258 669338 -5226 669574
rect -5846 609894 -5226 669338
rect -5846 609658 -5814 609894
rect -5578 609658 -5494 609894
rect -5258 609658 -5226 609894
rect -5846 609574 -5226 609658
rect -5846 609338 -5814 609574
rect -5578 609338 -5494 609574
rect -5258 609338 -5226 609574
rect -5846 549894 -5226 609338
rect -5846 549658 -5814 549894
rect -5578 549658 -5494 549894
rect -5258 549658 -5226 549894
rect -5846 549574 -5226 549658
rect -5846 549338 -5814 549574
rect -5578 549338 -5494 549574
rect -5258 549338 -5226 549574
rect -5846 489894 -5226 549338
rect -5846 489658 -5814 489894
rect -5578 489658 -5494 489894
rect -5258 489658 -5226 489894
rect -5846 489574 -5226 489658
rect -5846 489338 -5814 489574
rect -5578 489338 -5494 489574
rect -5258 489338 -5226 489574
rect -5846 429894 -5226 489338
rect -5846 429658 -5814 429894
rect -5578 429658 -5494 429894
rect -5258 429658 -5226 429894
rect -5846 429574 -5226 429658
rect -5846 429338 -5814 429574
rect -5578 429338 -5494 429574
rect -5258 429338 -5226 429574
rect -5846 369894 -5226 429338
rect -5846 369658 -5814 369894
rect -5578 369658 -5494 369894
rect -5258 369658 -5226 369894
rect -5846 369574 -5226 369658
rect -5846 369338 -5814 369574
rect -5578 369338 -5494 369574
rect -5258 369338 -5226 369574
rect -5846 309894 -5226 369338
rect -5846 309658 -5814 309894
rect -5578 309658 -5494 309894
rect -5258 309658 -5226 309894
rect -5846 309574 -5226 309658
rect -5846 309338 -5814 309574
rect -5578 309338 -5494 309574
rect -5258 309338 -5226 309574
rect -5846 249894 -5226 309338
rect -5846 249658 -5814 249894
rect -5578 249658 -5494 249894
rect -5258 249658 -5226 249894
rect -5846 249574 -5226 249658
rect -5846 249338 -5814 249574
rect -5578 249338 -5494 249574
rect -5258 249338 -5226 249574
rect -5846 189894 -5226 249338
rect -5846 189658 -5814 189894
rect -5578 189658 -5494 189894
rect -5258 189658 -5226 189894
rect -5846 189574 -5226 189658
rect -5846 189338 -5814 189574
rect -5578 189338 -5494 189574
rect -5258 189338 -5226 189574
rect -5846 129894 -5226 189338
rect -5846 129658 -5814 129894
rect -5578 129658 -5494 129894
rect -5258 129658 -5226 129894
rect -5846 129574 -5226 129658
rect -5846 129338 -5814 129574
rect -5578 129338 -5494 129574
rect -5258 129338 -5226 129574
rect -5846 69894 -5226 129338
rect -5846 69658 -5814 69894
rect -5578 69658 -5494 69894
rect -5258 69658 -5226 69894
rect -5846 69574 -5226 69658
rect -5846 69338 -5814 69574
rect -5578 69338 -5494 69574
rect -5258 69338 -5226 69574
rect -5846 9894 -5226 69338
rect -5846 9658 -5814 9894
rect -5578 9658 -5494 9894
rect -5258 9658 -5226 9894
rect -5846 9574 -5226 9658
rect -5846 9338 -5814 9574
rect -5578 9338 -5494 9574
rect -5258 9338 -5226 9574
rect -5846 -4186 -5226 9338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 696174 -4266 707162
rect -4886 695938 -4854 696174
rect -4618 695938 -4534 696174
rect -4298 695938 -4266 696174
rect -4886 695854 -4266 695938
rect -4886 695618 -4854 695854
rect -4618 695618 -4534 695854
rect -4298 695618 -4266 695854
rect -4886 636174 -4266 695618
rect -4886 635938 -4854 636174
rect -4618 635938 -4534 636174
rect -4298 635938 -4266 636174
rect -4886 635854 -4266 635938
rect -4886 635618 -4854 635854
rect -4618 635618 -4534 635854
rect -4298 635618 -4266 635854
rect -4886 576174 -4266 635618
rect -4886 575938 -4854 576174
rect -4618 575938 -4534 576174
rect -4298 575938 -4266 576174
rect -4886 575854 -4266 575938
rect -4886 575618 -4854 575854
rect -4618 575618 -4534 575854
rect -4298 575618 -4266 575854
rect -4886 516174 -4266 575618
rect -4886 515938 -4854 516174
rect -4618 515938 -4534 516174
rect -4298 515938 -4266 516174
rect -4886 515854 -4266 515938
rect -4886 515618 -4854 515854
rect -4618 515618 -4534 515854
rect -4298 515618 -4266 515854
rect -4886 456174 -4266 515618
rect -4886 455938 -4854 456174
rect -4618 455938 -4534 456174
rect -4298 455938 -4266 456174
rect -4886 455854 -4266 455938
rect -4886 455618 -4854 455854
rect -4618 455618 -4534 455854
rect -4298 455618 -4266 455854
rect -4886 396174 -4266 455618
rect -4886 395938 -4854 396174
rect -4618 395938 -4534 396174
rect -4298 395938 -4266 396174
rect -4886 395854 -4266 395938
rect -4886 395618 -4854 395854
rect -4618 395618 -4534 395854
rect -4298 395618 -4266 395854
rect -4886 336174 -4266 395618
rect -4886 335938 -4854 336174
rect -4618 335938 -4534 336174
rect -4298 335938 -4266 336174
rect -4886 335854 -4266 335938
rect -4886 335618 -4854 335854
rect -4618 335618 -4534 335854
rect -4298 335618 -4266 335854
rect -4886 276174 -4266 335618
rect -4886 275938 -4854 276174
rect -4618 275938 -4534 276174
rect -4298 275938 -4266 276174
rect -4886 275854 -4266 275938
rect -4886 275618 -4854 275854
rect -4618 275618 -4534 275854
rect -4298 275618 -4266 275854
rect -4886 216174 -4266 275618
rect -4886 215938 -4854 216174
rect -4618 215938 -4534 216174
rect -4298 215938 -4266 216174
rect -4886 215854 -4266 215938
rect -4886 215618 -4854 215854
rect -4618 215618 -4534 215854
rect -4298 215618 -4266 215854
rect -4886 156174 -4266 215618
rect -4886 155938 -4854 156174
rect -4618 155938 -4534 156174
rect -4298 155938 -4266 156174
rect -4886 155854 -4266 155938
rect -4886 155618 -4854 155854
rect -4618 155618 -4534 155854
rect -4298 155618 -4266 155854
rect -4886 96174 -4266 155618
rect -4886 95938 -4854 96174
rect -4618 95938 -4534 96174
rect -4298 95938 -4266 96174
rect -4886 95854 -4266 95938
rect -4886 95618 -4854 95854
rect -4618 95618 -4534 95854
rect -4298 95618 -4266 95854
rect -4886 36174 -4266 95618
rect -4886 35938 -4854 36174
rect -4618 35938 -4534 36174
rect -4298 35938 -4266 36174
rect -4886 35854 -4266 35938
rect -4886 35618 -4854 35854
rect -4618 35618 -4534 35854
rect -4298 35618 -4266 35854
rect -4886 -3226 -4266 35618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 666174 -3306 706202
rect 4514 706758 5134 707750
rect 4514 706522 4546 706758
rect 4782 706522 4866 706758
rect 5102 706522 5134 706758
rect 4514 706438 5134 706522
rect 4514 706202 4546 706438
rect 4782 706202 4866 706438
rect 5102 706202 5134 706438
rect -3926 665938 -3894 666174
rect -3658 665938 -3574 666174
rect -3338 665938 -3306 666174
rect -3926 665854 -3306 665938
rect -3926 665618 -3894 665854
rect -3658 665618 -3574 665854
rect -3338 665618 -3306 665854
rect -3926 606174 -3306 665618
rect -3926 605938 -3894 606174
rect -3658 605938 -3574 606174
rect -3338 605938 -3306 606174
rect -3926 605854 -3306 605938
rect -3926 605618 -3894 605854
rect -3658 605618 -3574 605854
rect -3338 605618 -3306 605854
rect -3926 546174 -3306 605618
rect -3926 545938 -3894 546174
rect -3658 545938 -3574 546174
rect -3338 545938 -3306 546174
rect -3926 545854 -3306 545938
rect -3926 545618 -3894 545854
rect -3658 545618 -3574 545854
rect -3338 545618 -3306 545854
rect -3926 486174 -3306 545618
rect -3926 485938 -3894 486174
rect -3658 485938 -3574 486174
rect -3338 485938 -3306 486174
rect -3926 485854 -3306 485938
rect -3926 485618 -3894 485854
rect -3658 485618 -3574 485854
rect -3338 485618 -3306 485854
rect -3926 426174 -3306 485618
rect -3926 425938 -3894 426174
rect -3658 425938 -3574 426174
rect -3338 425938 -3306 426174
rect -3926 425854 -3306 425938
rect -3926 425618 -3894 425854
rect -3658 425618 -3574 425854
rect -3338 425618 -3306 425854
rect -3926 366174 -3306 425618
rect -3926 365938 -3894 366174
rect -3658 365938 -3574 366174
rect -3338 365938 -3306 366174
rect -3926 365854 -3306 365938
rect -3926 365618 -3894 365854
rect -3658 365618 -3574 365854
rect -3338 365618 -3306 365854
rect -3926 306174 -3306 365618
rect -3926 305938 -3894 306174
rect -3658 305938 -3574 306174
rect -3338 305938 -3306 306174
rect -3926 305854 -3306 305938
rect -3926 305618 -3894 305854
rect -3658 305618 -3574 305854
rect -3338 305618 -3306 305854
rect -3926 246174 -3306 305618
rect -3926 245938 -3894 246174
rect -3658 245938 -3574 246174
rect -3338 245938 -3306 246174
rect -3926 245854 -3306 245938
rect -3926 245618 -3894 245854
rect -3658 245618 -3574 245854
rect -3338 245618 -3306 245854
rect -3926 186174 -3306 245618
rect -3926 185938 -3894 186174
rect -3658 185938 -3574 186174
rect -3338 185938 -3306 186174
rect -3926 185854 -3306 185938
rect -3926 185618 -3894 185854
rect -3658 185618 -3574 185854
rect -3338 185618 -3306 185854
rect -3926 126174 -3306 185618
rect -3926 125938 -3894 126174
rect -3658 125938 -3574 126174
rect -3338 125938 -3306 126174
rect -3926 125854 -3306 125938
rect -3926 125618 -3894 125854
rect -3658 125618 -3574 125854
rect -3338 125618 -3306 125854
rect -3926 66174 -3306 125618
rect -3926 65938 -3894 66174
rect -3658 65938 -3574 66174
rect -3338 65938 -3306 66174
rect -3926 65854 -3306 65938
rect -3926 65618 -3894 65854
rect -3658 65618 -3574 65854
rect -3338 65618 -3306 65854
rect -3926 6174 -3306 65618
rect -3926 5938 -3894 6174
rect -3658 5938 -3574 6174
rect -3338 5938 -3306 6174
rect -3926 5854 -3306 5938
rect -3926 5618 -3894 5854
rect -3658 5618 -3574 5854
rect -3338 5618 -3306 5854
rect -3926 -2266 -3306 5618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 692454 -2346 705242
rect -2966 692218 -2934 692454
rect -2698 692218 -2614 692454
rect -2378 692218 -2346 692454
rect -2966 692134 -2346 692218
rect -2966 691898 -2934 692134
rect -2698 691898 -2614 692134
rect -2378 691898 -2346 692134
rect -2966 632454 -2346 691898
rect -2966 632218 -2934 632454
rect -2698 632218 -2614 632454
rect -2378 632218 -2346 632454
rect -2966 632134 -2346 632218
rect -2966 631898 -2934 632134
rect -2698 631898 -2614 632134
rect -2378 631898 -2346 632134
rect -2966 572454 -2346 631898
rect -2966 572218 -2934 572454
rect -2698 572218 -2614 572454
rect -2378 572218 -2346 572454
rect -2966 572134 -2346 572218
rect -2966 571898 -2934 572134
rect -2698 571898 -2614 572134
rect -2378 571898 -2346 572134
rect -2966 512454 -2346 571898
rect -2966 512218 -2934 512454
rect -2698 512218 -2614 512454
rect -2378 512218 -2346 512454
rect -2966 512134 -2346 512218
rect -2966 511898 -2934 512134
rect -2698 511898 -2614 512134
rect -2378 511898 -2346 512134
rect -2966 452454 -2346 511898
rect -2966 452218 -2934 452454
rect -2698 452218 -2614 452454
rect -2378 452218 -2346 452454
rect -2966 452134 -2346 452218
rect -2966 451898 -2934 452134
rect -2698 451898 -2614 452134
rect -2378 451898 -2346 452134
rect -2966 392454 -2346 451898
rect -2966 392218 -2934 392454
rect -2698 392218 -2614 392454
rect -2378 392218 -2346 392454
rect -2966 392134 -2346 392218
rect -2966 391898 -2934 392134
rect -2698 391898 -2614 392134
rect -2378 391898 -2346 392134
rect -2966 332454 -2346 391898
rect -2966 332218 -2934 332454
rect -2698 332218 -2614 332454
rect -2378 332218 -2346 332454
rect -2966 332134 -2346 332218
rect -2966 331898 -2934 332134
rect -2698 331898 -2614 332134
rect -2378 331898 -2346 332134
rect -2966 272454 -2346 331898
rect -2966 272218 -2934 272454
rect -2698 272218 -2614 272454
rect -2378 272218 -2346 272454
rect -2966 272134 -2346 272218
rect -2966 271898 -2934 272134
rect -2698 271898 -2614 272134
rect -2378 271898 -2346 272134
rect -2966 212454 -2346 271898
rect -2966 212218 -2934 212454
rect -2698 212218 -2614 212454
rect -2378 212218 -2346 212454
rect -2966 212134 -2346 212218
rect -2966 211898 -2934 212134
rect -2698 211898 -2614 212134
rect -2378 211898 -2346 212134
rect -2966 152454 -2346 211898
rect -2966 152218 -2934 152454
rect -2698 152218 -2614 152454
rect -2378 152218 -2346 152454
rect -2966 152134 -2346 152218
rect -2966 151898 -2934 152134
rect -2698 151898 -2614 152134
rect -2378 151898 -2346 152134
rect -2966 92454 -2346 151898
rect -2966 92218 -2934 92454
rect -2698 92218 -2614 92454
rect -2378 92218 -2346 92454
rect -2966 92134 -2346 92218
rect -2966 91898 -2934 92134
rect -2698 91898 -2614 92134
rect -2378 91898 -2346 92134
rect -2966 32454 -2346 91898
rect -2966 32218 -2934 32454
rect -2698 32218 -2614 32454
rect -2378 32218 -2346 32454
rect -2966 32134 -2346 32218
rect -2966 31898 -2934 32134
rect -2698 31898 -2614 32134
rect -2378 31898 -2346 32134
rect -2966 -1306 -2346 31898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 662454 -1386 704282
rect -2006 662218 -1974 662454
rect -1738 662218 -1654 662454
rect -1418 662218 -1386 662454
rect -2006 662134 -1386 662218
rect -2006 661898 -1974 662134
rect -1738 661898 -1654 662134
rect -1418 661898 -1386 662134
rect -2006 602454 -1386 661898
rect -2006 602218 -1974 602454
rect -1738 602218 -1654 602454
rect -1418 602218 -1386 602454
rect -2006 602134 -1386 602218
rect -2006 601898 -1974 602134
rect -1738 601898 -1654 602134
rect -1418 601898 -1386 602134
rect -2006 542454 -1386 601898
rect -2006 542218 -1974 542454
rect -1738 542218 -1654 542454
rect -1418 542218 -1386 542454
rect -2006 542134 -1386 542218
rect -2006 541898 -1974 542134
rect -1738 541898 -1654 542134
rect -1418 541898 -1386 542134
rect -2006 482454 -1386 541898
rect -2006 482218 -1974 482454
rect -1738 482218 -1654 482454
rect -1418 482218 -1386 482454
rect -2006 482134 -1386 482218
rect -2006 481898 -1974 482134
rect -1738 481898 -1654 482134
rect -1418 481898 -1386 482134
rect -2006 422454 -1386 481898
rect -2006 422218 -1974 422454
rect -1738 422218 -1654 422454
rect -1418 422218 -1386 422454
rect -2006 422134 -1386 422218
rect -2006 421898 -1974 422134
rect -1738 421898 -1654 422134
rect -1418 421898 -1386 422134
rect -2006 362454 -1386 421898
rect -2006 362218 -1974 362454
rect -1738 362218 -1654 362454
rect -1418 362218 -1386 362454
rect -2006 362134 -1386 362218
rect -2006 361898 -1974 362134
rect -1738 361898 -1654 362134
rect -1418 361898 -1386 362134
rect -2006 302454 -1386 361898
rect -2006 302218 -1974 302454
rect -1738 302218 -1654 302454
rect -1418 302218 -1386 302454
rect -2006 302134 -1386 302218
rect -2006 301898 -1974 302134
rect -1738 301898 -1654 302134
rect -1418 301898 -1386 302134
rect -2006 242454 -1386 301898
rect -2006 242218 -1974 242454
rect -1738 242218 -1654 242454
rect -1418 242218 -1386 242454
rect -2006 242134 -1386 242218
rect -2006 241898 -1974 242134
rect -1738 241898 -1654 242134
rect -1418 241898 -1386 242134
rect -2006 182454 -1386 241898
rect -2006 182218 -1974 182454
rect -1738 182218 -1654 182454
rect -1418 182218 -1386 182454
rect -2006 182134 -1386 182218
rect -2006 181898 -1974 182134
rect -1738 181898 -1654 182134
rect -1418 181898 -1386 182134
rect -2006 122454 -1386 181898
rect -2006 122218 -1974 122454
rect -1738 122218 -1654 122454
rect -1418 122218 -1386 122454
rect -2006 122134 -1386 122218
rect -2006 121898 -1974 122134
rect -1738 121898 -1654 122134
rect -1418 121898 -1386 122134
rect -2006 62454 -1386 121898
rect -2006 62218 -1974 62454
rect -1738 62218 -1654 62454
rect -1418 62218 -1386 62454
rect -2006 62134 -1386 62218
rect -2006 61898 -1974 62134
rect -1738 61898 -1654 62134
rect -1418 61898 -1386 62134
rect -2006 2454 -1386 61898
rect -2006 2218 -1974 2454
rect -1738 2218 -1654 2454
rect -1418 2218 -1386 2454
rect -2006 2134 -1386 2218
rect -2006 1898 -1974 2134
rect -1738 1898 -1654 2134
rect -1418 1898 -1386 2134
rect -2006 -346 -1386 1898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 794 704838 1414 705830
rect 794 704602 826 704838
rect 1062 704602 1146 704838
rect 1382 704602 1414 704838
rect 794 704518 1414 704602
rect 794 704282 826 704518
rect 1062 704282 1146 704518
rect 1382 704282 1414 704518
rect 794 662454 1414 704282
rect 794 662218 826 662454
rect 1062 662218 1146 662454
rect 1382 662218 1414 662454
rect 794 662134 1414 662218
rect 794 661898 826 662134
rect 1062 661898 1146 662134
rect 1382 661898 1414 662134
rect 794 602454 1414 661898
rect 794 602218 826 602454
rect 1062 602218 1146 602454
rect 1382 602218 1414 602454
rect 794 602134 1414 602218
rect 794 601898 826 602134
rect 1062 601898 1146 602134
rect 1382 601898 1414 602134
rect 794 542454 1414 601898
rect 794 542218 826 542454
rect 1062 542218 1146 542454
rect 1382 542218 1414 542454
rect 794 542134 1414 542218
rect 794 541898 826 542134
rect 1062 541898 1146 542134
rect 1382 541898 1414 542134
rect 794 482454 1414 541898
rect 794 482218 826 482454
rect 1062 482218 1146 482454
rect 1382 482218 1414 482454
rect 794 482134 1414 482218
rect 794 481898 826 482134
rect 1062 481898 1146 482134
rect 1382 481898 1414 482134
rect 794 422454 1414 481898
rect 794 422218 826 422454
rect 1062 422218 1146 422454
rect 1382 422218 1414 422454
rect 794 422134 1414 422218
rect 794 421898 826 422134
rect 1062 421898 1146 422134
rect 1382 421898 1414 422134
rect 794 362454 1414 421898
rect 794 362218 826 362454
rect 1062 362218 1146 362454
rect 1382 362218 1414 362454
rect 794 362134 1414 362218
rect 794 361898 826 362134
rect 1062 361898 1146 362134
rect 1382 361898 1414 362134
rect 794 302454 1414 361898
rect 4514 666174 5134 706202
rect 4514 665938 4546 666174
rect 4782 665938 4866 666174
rect 5102 665938 5134 666174
rect 4514 665854 5134 665938
rect 4514 665618 4546 665854
rect 4782 665618 4866 665854
rect 5102 665618 5134 665854
rect 4514 606174 5134 665618
rect 4514 605938 4546 606174
rect 4782 605938 4866 606174
rect 5102 605938 5134 606174
rect 4514 605854 5134 605938
rect 4514 605618 4546 605854
rect 4782 605618 4866 605854
rect 5102 605618 5134 605854
rect 4514 546174 5134 605618
rect 4514 545938 4546 546174
rect 4782 545938 4866 546174
rect 5102 545938 5134 546174
rect 4514 545854 5134 545938
rect 4514 545618 4546 545854
rect 4782 545618 4866 545854
rect 5102 545618 5134 545854
rect 4514 486174 5134 545618
rect 4514 485938 4546 486174
rect 4782 485938 4866 486174
rect 5102 485938 5134 486174
rect 4514 485854 5134 485938
rect 4514 485618 4546 485854
rect 4782 485618 4866 485854
rect 5102 485618 5134 485854
rect 4514 426174 5134 485618
rect 4514 425938 4546 426174
rect 4782 425938 4866 426174
rect 5102 425938 5134 426174
rect 4514 425854 5134 425938
rect 4514 425618 4546 425854
rect 4782 425618 4866 425854
rect 5102 425618 5134 425854
rect 4514 366174 5134 425618
rect 4514 365938 4546 366174
rect 4782 365938 4866 366174
rect 5102 365938 5134 366174
rect 4514 365854 5134 365938
rect 4514 365618 4546 365854
rect 4782 365618 4866 365854
rect 5102 365618 5134 365854
rect 3371 358460 3437 358461
rect 3371 358396 3372 358460
rect 3436 358396 3437 358460
rect 3371 358395 3437 358396
rect 794 302218 826 302454
rect 1062 302218 1146 302454
rect 1382 302218 1414 302454
rect 794 302134 1414 302218
rect 794 301898 826 302134
rect 1062 301898 1146 302134
rect 1382 301898 1414 302134
rect 794 242454 1414 301898
rect 794 242218 826 242454
rect 1062 242218 1146 242454
rect 1382 242218 1414 242454
rect 794 242134 1414 242218
rect 794 241898 826 242134
rect 1062 241898 1146 242134
rect 1382 241898 1414 242134
rect 794 182454 1414 241898
rect 3374 204458 3434 358395
rect 4514 306174 5134 365618
rect 4514 305938 4546 306174
rect 4782 305938 4866 306174
rect 5102 305938 5134 306174
rect 4514 305854 5134 305938
rect 4514 305618 4546 305854
rect 4782 305618 4866 305854
rect 5102 305618 5134 305854
rect 4514 246174 5134 305618
rect 4514 245938 4546 246174
rect 4782 245938 4866 246174
rect 5102 245938 5134 246174
rect 4514 245854 5134 245938
rect 4514 245618 4546 245854
rect 4782 245618 4866 245854
rect 5102 245618 5134 245854
rect 794 182218 826 182454
rect 1062 182218 1146 182454
rect 1382 182218 1414 182454
rect 794 182134 1414 182218
rect 794 181898 826 182134
rect 1062 181898 1146 182134
rect 1382 181898 1414 182134
rect 794 122454 1414 181898
rect 794 122218 826 122454
rect 1062 122218 1146 122454
rect 1382 122218 1414 122454
rect 794 122134 1414 122218
rect 794 121898 826 122134
rect 1062 121898 1146 122134
rect 1382 121898 1414 122134
rect 794 62454 1414 121898
rect 794 62218 826 62454
rect 1062 62218 1146 62454
rect 1382 62218 1414 62454
rect 794 62134 1414 62218
rect 794 61898 826 62134
rect 1062 61898 1146 62134
rect 1382 61898 1414 62134
rect 794 2454 1414 61898
rect 794 2218 826 2454
rect 1062 2218 1146 2454
rect 1382 2218 1414 2454
rect 794 2134 1414 2218
rect 794 1898 826 2134
rect 1062 1898 1146 2134
rect 1382 1898 1414 2134
rect 794 -346 1414 1898
rect 794 -582 826 -346
rect 1062 -582 1146 -346
rect 1382 -582 1414 -346
rect 794 -666 1414 -582
rect 794 -902 826 -666
rect 1062 -902 1146 -666
rect 1382 -902 1414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 794 -1894 1414 -902
rect 4514 186174 5134 245618
rect 4514 185938 4546 186174
rect 4782 185938 4866 186174
rect 5102 185938 5134 186174
rect 4514 185854 5134 185938
rect 4514 185618 4546 185854
rect 4782 185618 4866 185854
rect 5102 185618 5134 185854
rect 4514 126174 5134 185618
rect 4514 125938 4546 126174
rect 4782 125938 4866 126174
rect 5102 125938 5134 126174
rect 4514 125854 5134 125938
rect 4514 125618 4546 125854
rect 4782 125618 4866 125854
rect 5102 125618 5134 125854
rect 4514 66174 5134 125618
rect 4514 65938 4546 66174
rect 4782 65938 4866 66174
rect 5102 65938 5134 66174
rect 4514 65854 5134 65938
rect 4514 65618 4546 65854
rect 4782 65618 4866 65854
rect 5102 65618 5134 65854
rect 4514 6174 5134 65618
rect 4514 5938 4546 6174
rect 4782 5938 4866 6174
rect 5102 5938 5134 6174
rect 4514 5854 5134 5938
rect 4514 5618 4546 5854
rect 4782 5618 4866 5854
rect 5102 5618 5134 5854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 4514 -2266 5134 5618
rect 4514 -2502 4546 -2266
rect 4782 -2502 4866 -2266
rect 5102 -2502 5134 -2266
rect 4514 -2586 5134 -2502
rect 4514 -2822 4546 -2586
rect 4782 -2822 4866 -2586
rect 5102 -2822 5134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 4514 -3814 5134 -2822
rect 8234 669894 8854 708122
rect 8234 669658 8266 669894
rect 8502 669658 8586 669894
rect 8822 669658 8854 669894
rect 8234 669574 8854 669658
rect 8234 669338 8266 669574
rect 8502 669338 8586 669574
rect 8822 669338 8854 669574
rect 8234 609894 8854 669338
rect 8234 609658 8266 609894
rect 8502 609658 8586 609894
rect 8822 609658 8854 609894
rect 8234 609574 8854 609658
rect 8234 609338 8266 609574
rect 8502 609338 8586 609574
rect 8822 609338 8854 609574
rect 8234 549894 8854 609338
rect 8234 549658 8266 549894
rect 8502 549658 8586 549894
rect 8822 549658 8854 549894
rect 8234 549574 8854 549658
rect 8234 549338 8266 549574
rect 8502 549338 8586 549574
rect 8822 549338 8854 549574
rect 8234 489894 8854 549338
rect 8234 489658 8266 489894
rect 8502 489658 8586 489894
rect 8822 489658 8854 489894
rect 8234 489574 8854 489658
rect 8234 489338 8266 489574
rect 8502 489338 8586 489574
rect 8822 489338 8854 489574
rect 8234 429894 8854 489338
rect 8234 429658 8266 429894
rect 8502 429658 8586 429894
rect 8822 429658 8854 429894
rect 8234 429574 8854 429658
rect 8234 429338 8266 429574
rect 8502 429338 8586 429574
rect 8822 429338 8854 429574
rect 8234 369894 8854 429338
rect 8234 369658 8266 369894
rect 8502 369658 8586 369894
rect 8822 369658 8854 369894
rect 8234 369574 8854 369658
rect 8234 369338 8266 369574
rect 8502 369338 8586 369574
rect 8822 369338 8854 369574
rect 8234 309894 8854 369338
rect 8234 309658 8266 309894
rect 8502 309658 8586 309894
rect 8822 309658 8854 309894
rect 8234 309574 8854 309658
rect 8234 309338 8266 309574
rect 8502 309338 8586 309574
rect 8822 309338 8854 309574
rect 8234 249894 8854 309338
rect 8234 249658 8266 249894
rect 8502 249658 8586 249894
rect 8822 249658 8854 249894
rect 8234 249574 8854 249658
rect 8234 249338 8266 249574
rect 8502 249338 8586 249574
rect 8822 249338 8854 249574
rect 8234 189894 8854 249338
rect 8234 189658 8266 189894
rect 8502 189658 8586 189894
rect 8822 189658 8854 189894
rect 8234 189574 8854 189658
rect 8234 189338 8266 189574
rect 8502 189338 8586 189574
rect 8822 189338 8854 189574
rect 8234 129894 8854 189338
rect 8234 129658 8266 129894
rect 8502 129658 8586 129894
rect 8822 129658 8854 129894
rect 8234 129574 8854 129658
rect 8234 129338 8266 129574
rect 8502 129338 8586 129574
rect 8822 129338 8854 129574
rect 8234 69894 8854 129338
rect 8234 69658 8266 69894
rect 8502 69658 8586 69894
rect 8822 69658 8854 69894
rect 8234 69574 8854 69658
rect 8234 69338 8266 69574
rect 8502 69338 8586 69574
rect 8822 69338 8854 69574
rect 8234 9894 8854 69338
rect 8234 9658 8266 9894
rect 8502 9658 8586 9894
rect 8822 9658 8854 9894
rect 8234 9574 8854 9658
rect 8234 9338 8266 9574
rect 8502 9338 8586 9574
rect 8822 9338 8854 9574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 8234 -4186 8854 9338
rect 8234 -4422 8266 -4186
rect 8502 -4422 8586 -4186
rect 8822 -4422 8854 -4186
rect 8234 -4506 8854 -4422
rect 8234 -4742 8266 -4506
rect 8502 -4742 8586 -4506
rect 8822 -4742 8854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 8234 -5734 8854 -4742
rect 11954 673614 12574 710042
rect 41954 711558 42574 711590
rect 41954 711322 41986 711558
rect 42222 711322 42306 711558
rect 42542 711322 42574 711558
rect 41954 711238 42574 711322
rect 41954 711002 41986 711238
rect 42222 711002 42306 711238
rect 42542 711002 42574 711238
rect 38234 709638 38854 709670
rect 38234 709402 38266 709638
rect 38502 709402 38586 709638
rect 38822 709402 38854 709638
rect 38234 709318 38854 709402
rect 38234 709082 38266 709318
rect 38502 709082 38586 709318
rect 38822 709082 38854 709318
rect 34514 707718 35134 707750
rect 34514 707482 34546 707718
rect 34782 707482 34866 707718
rect 35102 707482 35134 707718
rect 34514 707398 35134 707482
rect 34514 707162 34546 707398
rect 34782 707162 34866 707398
rect 35102 707162 35134 707398
rect 30794 705798 31414 705830
rect 30794 705562 30826 705798
rect 31062 705562 31146 705798
rect 31382 705562 31414 705798
rect 30794 705478 31414 705562
rect 30794 705242 30826 705478
rect 31062 705242 31146 705478
rect 31382 705242 31414 705478
rect 24715 699820 24781 699821
rect 24715 699756 24716 699820
rect 24780 699756 24781 699820
rect 24715 699755 24781 699756
rect 11954 673378 11986 673614
rect 12222 673378 12306 673614
rect 12542 673378 12574 673614
rect 11954 673294 12574 673378
rect 11954 673058 11986 673294
rect 12222 673058 12306 673294
rect 12542 673058 12574 673294
rect 11954 613614 12574 673058
rect 11954 613378 11986 613614
rect 12222 613378 12306 613614
rect 12542 613378 12574 613614
rect 11954 613294 12574 613378
rect 11954 613058 11986 613294
rect 12222 613058 12306 613294
rect 12542 613058 12574 613294
rect 11954 553614 12574 613058
rect 11954 553378 11986 553614
rect 12222 553378 12306 553614
rect 12542 553378 12574 553614
rect 11954 553294 12574 553378
rect 11954 553058 11986 553294
rect 12222 553058 12306 553294
rect 12542 553058 12574 553294
rect 11954 493614 12574 553058
rect 11954 493378 11986 493614
rect 12222 493378 12306 493614
rect 12542 493378 12574 493614
rect 11954 493294 12574 493378
rect 11954 493058 11986 493294
rect 12222 493058 12306 493294
rect 12542 493058 12574 493294
rect 11954 433614 12574 493058
rect 11954 433378 11986 433614
rect 12222 433378 12306 433614
rect 12542 433378 12574 433614
rect 11954 433294 12574 433378
rect 11954 433058 11986 433294
rect 12222 433058 12306 433294
rect 12542 433058 12574 433294
rect 11954 373614 12574 433058
rect 11954 373378 11986 373614
rect 12222 373378 12306 373614
rect 12542 373378 12574 373614
rect 11954 373294 12574 373378
rect 11954 373058 11986 373294
rect 12222 373058 12306 373294
rect 12542 373058 12574 373294
rect 11954 313614 12574 373058
rect 11954 313378 11986 313614
rect 12222 313378 12306 313614
rect 12542 313378 12574 313614
rect 11954 313294 12574 313378
rect 11954 313058 11986 313294
rect 12222 313058 12306 313294
rect 12542 313058 12574 313294
rect 11954 253614 12574 313058
rect 11954 253378 11986 253614
rect 12222 253378 12306 253614
rect 12542 253378 12574 253614
rect 11954 253294 12574 253378
rect 11954 253058 11986 253294
rect 12222 253058 12306 253294
rect 12542 253058 12574 253294
rect 11954 193614 12574 253058
rect 24718 247298 24778 699755
rect 30794 692454 31414 705242
rect 30794 692218 30826 692454
rect 31062 692218 31146 692454
rect 31382 692218 31414 692454
rect 30794 692134 31414 692218
rect 30794 691898 30826 692134
rect 31062 691898 31146 692134
rect 31382 691898 31414 692134
rect 30794 632454 31414 691898
rect 30794 632218 30826 632454
rect 31062 632218 31146 632454
rect 31382 632218 31414 632454
rect 30794 632134 31414 632218
rect 30794 631898 30826 632134
rect 31062 631898 31146 632134
rect 31382 631898 31414 632134
rect 30794 572454 31414 631898
rect 30794 572218 30826 572454
rect 31062 572218 31146 572454
rect 31382 572218 31414 572454
rect 30794 572134 31414 572218
rect 30794 571898 30826 572134
rect 31062 571898 31146 572134
rect 31382 571898 31414 572134
rect 30794 512454 31414 571898
rect 30794 512218 30826 512454
rect 31062 512218 31146 512454
rect 31382 512218 31414 512454
rect 30794 512134 31414 512218
rect 30794 511898 30826 512134
rect 31062 511898 31146 512134
rect 31382 511898 31414 512134
rect 30794 452454 31414 511898
rect 30794 452218 30826 452454
rect 31062 452218 31146 452454
rect 31382 452218 31414 452454
rect 30794 452134 31414 452218
rect 30794 451898 30826 452134
rect 31062 451898 31146 452134
rect 31382 451898 31414 452134
rect 30794 392454 31414 451898
rect 30794 392218 30826 392454
rect 31062 392218 31146 392454
rect 31382 392218 31414 392454
rect 30794 392134 31414 392218
rect 30794 391898 30826 392134
rect 31062 391898 31146 392134
rect 31382 391898 31414 392134
rect 30794 332454 31414 391898
rect 30794 332218 30826 332454
rect 31062 332218 31146 332454
rect 31382 332218 31414 332454
rect 30794 332134 31414 332218
rect 30794 331898 30826 332134
rect 31062 331898 31146 332134
rect 31382 331898 31414 332134
rect 30794 272454 31414 331898
rect 30794 272218 30826 272454
rect 31062 272218 31146 272454
rect 31382 272218 31414 272454
rect 30794 272134 31414 272218
rect 30794 271898 30826 272134
rect 31062 271898 31146 272134
rect 31382 271898 31414 272134
rect 11954 193378 11986 193614
rect 12222 193378 12306 193614
rect 12542 193378 12574 193614
rect 11954 193294 12574 193378
rect 11954 193058 11986 193294
rect 12222 193058 12306 193294
rect 12542 193058 12574 193294
rect 11954 133614 12574 193058
rect 11954 133378 11986 133614
rect 12222 133378 12306 133614
rect 12542 133378 12574 133614
rect 11954 133294 12574 133378
rect 11954 133058 11986 133294
rect 12222 133058 12306 133294
rect 12542 133058 12574 133294
rect 11954 73614 12574 133058
rect 11954 73378 11986 73614
rect 12222 73378 12306 73614
rect 12542 73378 12574 73614
rect 11954 73294 12574 73378
rect 11954 73058 11986 73294
rect 12222 73058 12306 73294
rect 12542 73058 12574 73294
rect 11954 13614 12574 73058
rect 11954 13378 11986 13614
rect 12222 13378 12306 13614
rect 12542 13378 12574 13614
rect 11954 13294 12574 13378
rect 11954 13058 11986 13294
rect 12222 13058 12306 13294
rect 12542 13058 12574 13294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 11954 -6106 12574 13058
rect 30794 212454 31414 271898
rect 30794 212218 30826 212454
rect 31062 212218 31146 212454
rect 31382 212218 31414 212454
rect 30794 212134 31414 212218
rect 30794 211898 30826 212134
rect 31062 211898 31146 212134
rect 31382 211898 31414 212134
rect 30794 152454 31414 211898
rect 30794 152218 30826 152454
rect 31062 152218 31146 152454
rect 31382 152218 31414 152454
rect 30794 152134 31414 152218
rect 30794 151898 30826 152134
rect 31062 151898 31146 152134
rect 31382 151898 31414 152134
rect 30794 92454 31414 151898
rect 30794 92218 30826 92454
rect 31062 92218 31146 92454
rect 31382 92218 31414 92454
rect 30794 92134 31414 92218
rect 30794 91898 30826 92134
rect 31062 91898 31146 92134
rect 31382 91898 31414 92134
rect 30794 32454 31414 91898
rect 30794 32218 30826 32454
rect 31062 32218 31146 32454
rect 31382 32218 31414 32454
rect 30794 32134 31414 32218
rect 30794 31898 30826 32134
rect 31062 31898 31146 32134
rect 31382 31898 31414 32134
rect 30794 -1306 31414 31898
rect 30794 -1542 30826 -1306
rect 31062 -1542 31146 -1306
rect 31382 -1542 31414 -1306
rect 30794 -1626 31414 -1542
rect 30794 -1862 30826 -1626
rect 31062 -1862 31146 -1626
rect 31382 -1862 31414 -1626
rect 30794 -1894 31414 -1862
rect 34514 696174 35134 707162
rect 34514 695938 34546 696174
rect 34782 695938 34866 696174
rect 35102 695938 35134 696174
rect 34514 695854 35134 695938
rect 34514 695618 34546 695854
rect 34782 695618 34866 695854
rect 35102 695618 35134 695854
rect 34514 636174 35134 695618
rect 34514 635938 34546 636174
rect 34782 635938 34866 636174
rect 35102 635938 35134 636174
rect 34514 635854 35134 635938
rect 34514 635618 34546 635854
rect 34782 635618 34866 635854
rect 35102 635618 35134 635854
rect 34514 576174 35134 635618
rect 34514 575938 34546 576174
rect 34782 575938 34866 576174
rect 35102 575938 35134 576174
rect 34514 575854 35134 575938
rect 34514 575618 34546 575854
rect 34782 575618 34866 575854
rect 35102 575618 35134 575854
rect 34514 516174 35134 575618
rect 34514 515938 34546 516174
rect 34782 515938 34866 516174
rect 35102 515938 35134 516174
rect 34514 515854 35134 515938
rect 34514 515618 34546 515854
rect 34782 515618 34866 515854
rect 35102 515618 35134 515854
rect 34514 456174 35134 515618
rect 34514 455938 34546 456174
rect 34782 455938 34866 456174
rect 35102 455938 35134 456174
rect 34514 455854 35134 455938
rect 34514 455618 34546 455854
rect 34782 455618 34866 455854
rect 35102 455618 35134 455854
rect 34514 396174 35134 455618
rect 34514 395938 34546 396174
rect 34782 395938 34866 396174
rect 35102 395938 35134 396174
rect 34514 395854 35134 395938
rect 34514 395618 34546 395854
rect 34782 395618 34866 395854
rect 35102 395618 35134 395854
rect 34514 336174 35134 395618
rect 34514 335938 34546 336174
rect 34782 335938 34866 336174
rect 35102 335938 35134 336174
rect 34514 335854 35134 335938
rect 34514 335618 34546 335854
rect 34782 335618 34866 335854
rect 35102 335618 35134 335854
rect 34514 276174 35134 335618
rect 34514 275938 34546 276174
rect 34782 275938 34866 276174
rect 35102 275938 35134 276174
rect 34514 275854 35134 275938
rect 34514 275618 34546 275854
rect 34782 275618 34866 275854
rect 35102 275618 35134 275854
rect 34514 216174 35134 275618
rect 34514 215938 34546 216174
rect 34782 215938 34866 216174
rect 35102 215938 35134 216174
rect 34514 215854 35134 215938
rect 34514 215618 34546 215854
rect 34782 215618 34866 215854
rect 35102 215618 35134 215854
rect 34514 156174 35134 215618
rect 34514 155938 34546 156174
rect 34782 155938 34866 156174
rect 35102 155938 35134 156174
rect 34514 155854 35134 155938
rect 34514 155618 34546 155854
rect 34782 155618 34866 155854
rect 35102 155618 35134 155854
rect 34514 96174 35134 155618
rect 34514 95938 34546 96174
rect 34782 95938 34866 96174
rect 35102 95938 35134 96174
rect 34514 95854 35134 95938
rect 34514 95618 34546 95854
rect 34782 95618 34866 95854
rect 35102 95618 35134 95854
rect 34514 36174 35134 95618
rect 34514 35938 34546 36174
rect 34782 35938 34866 36174
rect 35102 35938 35134 36174
rect 34514 35854 35134 35938
rect 34514 35618 34546 35854
rect 34782 35618 34866 35854
rect 35102 35618 35134 35854
rect 34514 -3226 35134 35618
rect 34514 -3462 34546 -3226
rect 34782 -3462 34866 -3226
rect 35102 -3462 35134 -3226
rect 34514 -3546 35134 -3462
rect 34514 -3782 34546 -3546
rect 34782 -3782 34866 -3546
rect 35102 -3782 35134 -3546
rect 34514 -3814 35134 -3782
rect 38234 699894 38854 709082
rect 38234 699658 38266 699894
rect 38502 699658 38586 699894
rect 38822 699658 38854 699894
rect 38234 699574 38854 699658
rect 38234 699338 38266 699574
rect 38502 699338 38586 699574
rect 38822 699338 38854 699574
rect 38234 639894 38854 699338
rect 38234 639658 38266 639894
rect 38502 639658 38586 639894
rect 38822 639658 38854 639894
rect 38234 639574 38854 639658
rect 38234 639338 38266 639574
rect 38502 639338 38586 639574
rect 38822 639338 38854 639574
rect 38234 579894 38854 639338
rect 38234 579658 38266 579894
rect 38502 579658 38586 579894
rect 38822 579658 38854 579894
rect 38234 579574 38854 579658
rect 38234 579338 38266 579574
rect 38502 579338 38586 579574
rect 38822 579338 38854 579574
rect 38234 519894 38854 579338
rect 38234 519658 38266 519894
rect 38502 519658 38586 519894
rect 38822 519658 38854 519894
rect 38234 519574 38854 519658
rect 38234 519338 38266 519574
rect 38502 519338 38586 519574
rect 38822 519338 38854 519574
rect 38234 459894 38854 519338
rect 38234 459658 38266 459894
rect 38502 459658 38586 459894
rect 38822 459658 38854 459894
rect 38234 459574 38854 459658
rect 38234 459338 38266 459574
rect 38502 459338 38586 459574
rect 38822 459338 38854 459574
rect 38234 399894 38854 459338
rect 38234 399658 38266 399894
rect 38502 399658 38586 399894
rect 38822 399658 38854 399894
rect 38234 399574 38854 399658
rect 38234 399338 38266 399574
rect 38502 399338 38586 399574
rect 38822 399338 38854 399574
rect 38234 339894 38854 399338
rect 38234 339658 38266 339894
rect 38502 339658 38586 339894
rect 38822 339658 38854 339894
rect 38234 339574 38854 339658
rect 38234 339338 38266 339574
rect 38502 339338 38586 339574
rect 38822 339338 38854 339574
rect 38234 279894 38854 339338
rect 38234 279658 38266 279894
rect 38502 279658 38586 279894
rect 38822 279658 38854 279894
rect 38234 279574 38854 279658
rect 38234 279338 38266 279574
rect 38502 279338 38586 279574
rect 38822 279338 38854 279574
rect 38234 219894 38854 279338
rect 38234 219658 38266 219894
rect 38502 219658 38586 219894
rect 38822 219658 38854 219894
rect 38234 219574 38854 219658
rect 38234 219338 38266 219574
rect 38502 219338 38586 219574
rect 38822 219338 38854 219574
rect 38234 159894 38854 219338
rect 38234 159658 38266 159894
rect 38502 159658 38586 159894
rect 38822 159658 38854 159894
rect 38234 159574 38854 159658
rect 38234 159338 38266 159574
rect 38502 159338 38586 159574
rect 38822 159338 38854 159574
rect 38234 99894 38854 159338
rect 38234 99658 38266 99894
rect 38502 99658 38586 99894
rect 38822 99658 38854 99894
rect 38234 99574 38854 99658
rect 38234 99338 38266 99574
rect 38502 99338 38586 99574
rect 38822 99338 38854 99574
rect 38234 39894 38854 99338
rect 38234 39658 38266 39894
rect 38502 39658 38586 39894
rect 38822 39658 38854 39894
rect 38234 39574 38854 39658
rect 38234 39338 38266 39574
rect 38502 39338 38586 39574
rect 38822 39338 38854 39574
rect 38234 -5146 38854 39338
rect 38234 -5382 38266 -5146
rect 38502 -5382 38586 -5146
rect 38822 -5382 38854 -5146
rect 38234 -5466 38854 -5382
rect 38234 -5702 38266 -5466
rect 38502 -5702 38586 -5466
rect 38822 -5702 38854 -5466
rect 38234 -5734 38854 -5702
rect 41954 643614 42574 711002
rect 71954 710598 72574 711590
rect 71954 710362 71986 710598
rect 72222 710362 72306 710598
rect 72542 710362 72574 710598
rect 71954 710278 72574 710362
rect 71954 710042 71986 710278
rect 72222 710042 72306 710278
rect 72542 710042 72574 710278
rect 68234 708678 68854 709670
rect 68234 708442 68266 708678
rect 68502 708442 68586 708678
rect 68822 708442 68854 708678
rect 68234 708358 68854 708442
rect 68234 708122 68266 708358
rect 68502 708122 68586 708358
rect 68822 708122 68854 708358
rect 64514 706758 65134 707750
rect 64514 706522 64546 706758
rect 64782 706522 64866 706758
rect 65102 706522 65134 706758
rect 64514 706438 65134 706522
rect 64514 706202 64546 706438
rect 64782 706202 64866 706438
rect 65102 706202 65134 706438
rect 41954 643378 41986 643614
rect 42222 643378 42306 643614
rect 42542 643378 42574 643614
rect 41954 643294 42574 643378
rect 41954 643058 41986 643294
rect 42222 643058 42306 643294
rect 42542 643058 42574 643294
rect 41954 583614 42574 643058
rect 41954 583378 41986 583614
rect 42222 583378 42306 583614
rect 42542 583378 42574 583614
rect 41954 583294 42574 583378
rect 41954 583058 41986 583294
rect 42222 583058 42306 583294
rect 42542 583058 42574 583294
rect 41954 523614 42574 583058
rect 41954 523378 41986 523614
rect 42222 523378 42306 523614
rect 42542 523378 42574 523614
rect 41954 523294 42574 523378
rect 41954 523058 41986 523294
rect 42222 523058 42306 523294
rect 42542 523058 42574 523294
rect 41954 463614 42574 523058
rect 41954 463378 41986 463614
rect 42222 463378 42306 463614
rect 42542 463378 42574 463614
rect 41954 463294 42574 463378
rect 41954 463058 41986 463294
rect 42222 463058 42306 463294
rect 42542 463058 42574 463294
rect 41954 403614 42574 463058
rect 41954 403378 41986 403614
rect 42222 403378 42306 403614
rect 42542 403378 42574 403614
rect 41954 403294 42574 403378
rect 41954 403058 41986 403294
rect 42222 403058 42306 403294
rect 42542 403058 42574 403294
rect 41954 343614 42574 403058
rect 41954 343378 41986 343614
rect 42222 343378 42306 343614
rect 42542 343378 42574 343614
rect 41954 343294 42574 343378
rect 41954 343058 41986 343294
rect 42222 343058 42306 343294
rect 42542 343058 42574 343294
rect 41954 283614 42574 343058
rect 41954 283378 41986 283614
rect 42222 283378 42306 283614
rect 42542 283378 42574 283614
rect 41954 283294 42574 283378
rect 41954 283058 41986 283294
rect 42222 283058 42306 283294
rect 42542 283058 42574 283294
rect 41954 223614 42574 283058
rect 41954 223378 41986 223614
rect 42222 223378 42306 223614
rect 42542 223378 42574 223614
rect 41954 223294 42574 223378
rect 41954 223058 41986 223294
rect 42222 223058 42306 223294
rect 42542 223058 42574 223294
rect 41954 163614 42574 223058
rect 41954 163378 41986 163614
rect 42222 163378 42306 163614
rect 42542 163378 42574 163614
rect 41954 163294 42574 163378
rect 41954 163058 41986 163294
rect 42222 163058 42306 163294
rect 42542 163058 42574 163294
rect 41954 103614 42574 163058
rect 41954 103378 41986 103614
rect 42222 103378 42306 103614
rect 42542 103378 42574 103614
rect 41954 103294 42574 103378
rect 41954 103058 41986 103294
rect 42222 103058 42306 103294
rect 42542 103058 42574 103294
rect 41954 43614 42574 103058
rect 41954 43378 41986 43614
rect 42222 43378 42306 43614
rect 42542 43378 42574 43614
rect 41954 43294 42574 43378
rect 41954 43058 41986 43294
rect 42222 43058 42306 43294
rect 42542 43058 42574 43294
rect 11954 -6342 11986 -6106
rect 12222 -6342 12306 -6106
rect 12542 -6342 12574 -6106
rect 11954 -6426 12574 -6342
rect 11954 -6662 11986 -6426
rect 12222 -6662 12306 -6426
rect 12542 -6662 12574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 11954 -7654 12574 -6662
rect 41954 -7066 42574 43058
rect 60794 704838 61414 705830
rect 60794 704602 60826 704838
rect 61062 704602 61146 704838
rect 61382 704602 61414 704838
rect 60794 704518 61414 704602
rect 60794 704282 60826 704518
rect 61062 704282 61146 704518
rect 61382 704282 61414 704518
rect 60794 662454 61414 704282
rect 60794 662218 60826 662454
rect 61062 662218 61146 662454
rect 61382 662218 61414 662454
rect 60794 662134 61414 662218
rect 60794 661898 60826 662134
rect 61062 661898 61146 662134
rect 61382 661898 61414 662134
rect 60794 602454 61414 661898
rect 60794 602218 60826 602454
rect 61062 602218 61146 602454
rect 61382 602218 61414 602454
rect 60794 602134 61414 602218
rect 60794 601898 60826 602134
rect 61062 601898 61146 602134
rect 61382 601898 61414 602134
rect 60794 542454 61414 601898
rect 60794 542218 60826 542454
rect 61062 542218 61146 542454
rect 61382 542218 61414 542454
rect 60794 542134 61414 542218
rect 60794 541898 60826 542134
rect 61062 541898 61146 542134
rect 61382 541898 61414 542134
rect 60794 482454 61414 541898
rect 60794 482218 60826 482454
rect 61062 482218 61146 482454
rect 61382 482218 61414 482454
rect 60794 482134 61414 482218
rect 60794 481898 60826 482134
rect 61062 481898 61146 482134
rect 61382 481898 61414 482134
rect 60794 422454 61414 481898
rect 60794 422218 60826 422454
rect 61062 422218 61146 422454
rect 61382 422218 61414 422454
rect 60794 422134 61414 422218
rect 60794 421898 60826 422134
rect 61062 421898 61146 422134
rect 61382 421898 61414 422134
rect 60794 362454 61414 421898
rect 60794 362218 60826 362454
rect 61062 362218 61146 362454
rect 61382 362218 61414 362454
rect 60794 362134 61414 362218
rect 60794 361898 60826 362134
rect 61062 361898 61146 362134
rect 61382 361898 61414 362134
rect 60794 302454 61414 361898
rect 60794 302218 60826 302454
rect 61062 302218 61146 302454
rect 61382 302218 61414 302454
rect 60794 302134 61414 302218
rect 60794 301898 60826 302134
rect 61062 301898 61146 302134
rect 61382 301898 61414 302134
rect 60794 242454 61414 301898
rect 60794 242218 60826 242454
rect 61062 242218 61146 242454
rect 61382 242218 61414 242454
rect 60794 242134 61414 242218
rect 60794 241898 60826 242134
rect 61062 241898 61146 242134
rect 61382 241898 61414 242134
rect 60794 182454 61414 241898
rect 60794 182218 60826 182454
rect 61062 182218 61146 182454
rect 61382 182218 61414 182454
rect 60794 182134 61414 182218
rect 60794 181898 60826 182134
rect 61062 181898 61146 182134
rect 61382 181898 61414 182134
rect 60794 122454 61414 181898
rect 60794 122218 60826 122454
rect 61062 122218 61146 122454
rect 61382 122218 61414 122454
rect 60794 122134 61414 122218
rect 60794 121898 60826 122134
rect 61062 121898 61146 122134
rect 61382 121898 61414 122134
rect 60794 62454 61414 121898
rect 60794 62218 60826 62454
rect 61062 62218 61146 62454
rect 61382 62218 61414 62454
rect 60794 62134 61414 62218
rect 60794 61898 60826 62134
rect 61062 61898 61146 62134
rect 61382 61898 61414 62134
rect 60794 2454 61414 61898
rect 60794 2218 60826 2454
rect 61062 2218 61146 2454
rect 61382 2218 61414 2454
rect 60794 2134 61414 2218
rect 60794 1898 60826 2134
rect 61062 1898 61146 2134
rect 61382 1898 61414 2134
rect 60794 -346 61414 1898
rect 60794 -582 60826 -346
rect 61062 -582 61146 -346
rect 61382 -582 61414 -346
rect 60794 -666 61414 -582
rect 60794 -902 60826 -666
rect 61062 -902 61146 -666
rect 61382 -902 61414 -666
rect 60794 -1894 61414 -902
rect 64514 666174 65134 706202
rect 64514 665938 64546 666174
rect 64782 665938 64866 666174
rect 65102 665938 65134 666174
rect 64514 665854 65134 665938
rect 64514 665618 64546 665854
rect 64782 665618 64866 665854
rect 65102 665618 65134 665854
rect 64514 606174 65134 665618
rect 64514 605938 64546 606174
rect 64782 605938 64866 606174
rect 65102 605938 65134 606174
rect 64514 605854 65134 605938
rect 64514 605618 64546 605854
rect 64782 605618 64866 605854
rect 65102 605618 65134 605854
rect 64514 546174 65134 605618
rect 64514 545938 64546 546174
rect 64782 545938 64866 546174
rect 65102 545938 65134 546174
rect 64514 545854 65134 545938
rect 64514 545618 64546 545854
rect 64782 545618 64866 545854
rect 65102 545618 65134 545854
rect 64514 486174 65134 545618
rect 64514 485938 64546 486174
rect 64782 485938 64866 486174
rect 65102 485938 65134 486174
rect 64514 485854 65134 485938
rect 64514 485618 64546 485854
rect 64782 485618 64866 485854
rect 65102 485618 65134 485854
rect 64514 426174 65134 485618
rect 64514 425938 64546 426174
rect 64782 425938 64866 426174
rect 65102 425938 65134 426174
rect 64514 425854 65134 425938
rect 64514 425618 64546 425854
rect 64782 425618 64866 425854
rect 65102 425618 65134 425854
rect 64514 366174 65134 425618
rect 64514 365938 64546 366174
rect 64782 365938 64866 366174
rect 65102 365938 65134 366174
rect 64514 365854 65134 365938
rect 64514 365618 64546 365854
rect 64782 365618 64866 365854
rect 65102 365618 65134 365854
rect 64514 306174 65134 365618
rect 64514 305938 64546 306174
rect 64782 305938 64866 306174
rect 65102 305938 65134 306174
rect 64514 305854 65134 305938
rect 64514 305618 64546 305854
rect 64782 305618 64866 305854
rect 65102 305618 65134 305854
rect 64514 246174 65134 305618
rect 64514 245938 64546 246174
rect 64782 245938 64866 246174
rect 65102 245938 65134 246174
rect 64514 245854 65134 245938
rect 64514 245618 64546 245854
rect 64782 245618 64866 245854
rect 65102 245618 65134 245854
rect 64514 186174 65134 245618
rect 64514 185938 64546 186174
rect 64782 185938 64866 186174
rect 65102 185938 65134 186174
rect 64514 185854 65134 185938
rect 64514 185618 64546 185854
rect 64782 185618 64866 185854
rect 65102 185618 65134 185854
rect 64514 126174 65134 185618
rect 64514 125938 64546 126174
rect 64782 125938 64866 126174
rect 65102 125938 65134 126174
rect 64514 125854 65134 125938
rect 64514 125618 64546 125854
rect 64782 125618 64866 125854
rect 65102 125618 65134 125854
rect 64514 66174 65134 125618
rect 64514 65938 64546 66174
rect 64782 65938 64866 66174
rect 65102 65938 65134 66174
rect 64514 65854 65134 65938
rect 64514 65618 64546 65854
rect 64782 65618 64866 65854
rect 65102 65618 65134 65854
rect 64514 6174 65134 65618
rect 64514 5938 64546 6174
rect 64782 5938 64866 6174
rect 65102 5938 65134 6174
rect 64514 5854 65134 5938
rect 64514 5618 64546 5854
rect 64782 5618 64866 5854
rect 65102 5618 65134 5854
rect 64514 -2266 65134 5618
rect 64514 -2502 64546 -2266
rect 64782 -2502 64866 -2266
rect 65102 -2502 65134 -2266
rect 64514 -2586 65134 -2502
rect 64514 -2822 64546 -2586
rect 64782 -2822 64866 -2586
rect 65102 -2822 65134 -2586
rect 64514 -3814 65134 -2822
rect 68234 669894 68854 708122
rect 68234 669658 68266 669894
rect 68502 669658 68586 669894
rect 68822 669658 68854 669894
rect 68234 669574 68854 669658
rect 68234 669338 68266 669574
rect 68502 669338 68586 669574
rect 68822 669338 68854 669574
rect 68234 609894 68854 669338
rect 68234 609658 68266 609894
rect 68502 609658 68586 609894
rect 68822 609658 68854 609894
rect 68234 609574 68854 609658
rect 68234 609338 68266 609574
rect 68502 609338 68586 609574
rect 68822 609338 68854 609574
rect 68234 549894 68854 609338
rect 68234 549658 68266 549894
rect 68502 549658 68586 549894
rect 68822 549658 68854 549894
rect 68234 549574 68854 549658
rect 68234 549338 68266 549574
rect 68502 549338 68586 549574
rect 68822 549338 68854 549574
rect 68234 489894 68854 549338
rect 68234 489658 68266 489894
rect 68502 489658 68586 489894
rect 68822 489658 68854 489894
rect 68234 489574 68854 489658
rect 68234 489338 68266 489574
rect 68502 489338 68586 489574
rect 68822 489338 68854 489574
rect 68234 429894 68854 489338
rect 68234 429658 68266 429894
rect 68502 429658 68586 429894
rect 68822 429658 68854 429894
rect 68234 429574 68854 429658
rect 68234 429338 68266 429574
rect 68502 429338 68586 429574
rect 68822 429338 68854 429574
rect 68234 369894 68854 429338
rect 68234 369658 68266 369894
rect 68502 369658 68586 369894
rect 68822 369658 68854 369894
rect 68234 369574 68854 369658
rect 68234 369338 68266 369574
rect 68502 369338 68586 369574
rect 68822 369338 68854 369574
rect 68234 309894 68854 369338
rect 68234 309658 68266 309894
rect 68502 309658 68586 309894
rect 68822 309658 68854 309894
rect 68234 309574 68854 309658
rect 68234 309338 68266 309574
rect 68502 309338 68586 309574
rect 68822 309338 68854 309574
rect 68234 249894 68854 309338
rect 68234 249658 68266 249894
rect 68502 249658 68586 249894
rect 68822 249658 68854 249894
rect 68234 249574 68854 249658
rect 68234 249338 68266 249574
rect 68502 249338 68586 249574
rect 68822 249338 68854 249574
rect 68234 189894 68854 249338
rect 68234 189658 68266 189894
rect 68502 189658 68586 189894
rect 68822 189658 68854 189894
rect 68234 189574 68854 189658
rect 68234 189338 68266 189574
rect 68502 189338 68586 189574
rect 68822 189338 68854 189574
rect 68234 129894 68854 189338
rect 68234 129658 68266 129894
rect 68502 129658 68586 129894
rect 68822 129658 68854 129894
rect 68234 129574 68854 129658
rect 68234 129338 68266 129574
rect 68502 129338 68586 129574
rect 68822 129338 68854 129574
rect 68234 69894 68854 129338
rect 68234 69658 68266 69894
rect 68502 69658 68586 69894
rect 68822 69658 68854 69894
rect 68234 69574 68854 69658
rect 68234 69338 68266 69574
rect 68502 69338 68586 69574
rect 68822 69338 68854 69574
rect 68234 9894 68854 69338
rect 68234 9658 68266 9894
rect 68502 9658 68586 9894
rect 68822 9658 68854 9894
rect 68234 9574 68854 9658
rect 68234 9338 68266 9574
rect 68502 9338 68586 9574
rect 68822 9338 68854 9574
rect 68234 -4186 68854 9338
rect 68234 -4422 68266 -4186
rect 68502 -4422 68586 -4186
rect 68822 -4422 68854 -4186
rect 68234 -4506 68854 -4422
rect 68234 -4742 68266 -4506
rect 68502 -4742 68586 -4506
rect 68822 -4742 68854 -4506
rect 68234 -5734 68854 -4742
rect 71954 673614 72574 710042
rect 101954 711558 102574 711590
rect 101954 711322 101986 711558
rect 102222 711322 102306 711558
rect 102542 711322 102574 711558
rect 101954 711238 102574 711322
rect 101954 711002 101986 711238
rect 102222 711002 102306 711238
rect 102542 711002 102574 711238
rect 98234 709638 98854 709670
rect 98234 709402 98266 709638
rect 98502 709402 98586 709638
rect 98822 709402 98854 709638
rect 98234 709318 98854 709402
rect 98234 709082 98266 709318
rect 98502 709082 98586 709318
rect 98822 709082 98854 709318
rect 94514 707718 95134 707750
rect 94514 707482 94546 707718
rect 94782 707482 94866 707718
rect 95102 707482 95134 707718
rect 94514 707398 95134 707482
rect 94514 707162 94546 707398
rect 94782 707162 94866 707398
rect 95102 707162 95134 707398
rect 71954 673378 71986 673614
rect 72222 673378 72306 673614
rect 72542 673378 72574 673614
rect 71954 673294 72574 673378
rect 71954 673058 71986 673294
rect 72222 673058 72306 673294
rect 72542 673058 72574 673294
rect 71954 613614 72574 673058
rect 71954 613378 71986 613614
rect 72222 613378 72306 613614
rect 72542 613378 72574 613614
rect 71954 613294 72574 613378
rect 71954 613058 71986 613294
rect 72222 613058 72306 613294
rect 72542 613058 72574 613294
rect 71954 553614 72574 613058
rect 71954 553378 71986 553614
rect 72222 553378 72306 553614
rect 72542 553378 72574 553614
rect 71954 553294 72574 553378
rect 71954 553058 71986 553294
rect 72222 553058 72306 553294
rect 72542 553058 72574 553294
rect 71954 493614 72574 553058
rect 71954 493378 71986 493614
rect 72222 493378 72306 493614
rect 72542 493378 72574 493614
rect 71954 493294 72574 493378
rect 71954 493058 71986 493294
rect 72222 493058 72306 493294
rect 72542 493058 72574 493294
rect 71954 433614 72574 493058
rect 71954 433378 71986 433614
rect 72222 433378 72306 433614
rect 72542 433378 72574 433614
rect 71954 433294 72574 433378
rect 71954 433058 71986 433294
rect 72222 433058 72306 433294
rect 72542 433058 72574 433294
rect 71954 373614 72574 433058
rect 71954 373378 71986 373614
rect 72222 373378 72306 373614
rect 72542 373378 72574 373614
rect 71954 373294 72574 373378
rect 71954 373058 71986 373294
rect 72222 373058 72306 373294
rect 72542 373058 72574 373294
rect 71954 313614 72574 373058
rect 71954 313378 71986 313614
rect 72222 313378 72306 313614
rect 72542 313378 72574 313614
rect 71954 313294 72574 313378
rect 71954 313058 71986 313294
rect 72222 313058 72306 313294
rect 72542 313058 72574 313294
rect 71954 253614 72574 313058
rect 71954 253378 71986 253614
rect 72222 253378 72306 253614
rect 72542 253378 72574 253614
rect 71954 253294 72574 253378
rect 71954 253058 71986 253294
rect 72222 253058 72306 253294
rect 72542 253058 72574 253294
rect 71954 193614 72574 253058
rect 71954 193378 71986 193614
rect 72222 193378 72306 193614
rect 72542 193378 72574 193614
rect 71954 193294 72574 193378
rect 71954 193058 71986 193294
rect 72222 193058 72306 193294
rect 72542 193058 72574 193294
rect 71954 133614 72574 193058
rect 71954 133378 71986 133614
rect 72222 133378 72306 133614
rect 72542 133378 72574 133614
rect 71954 133294 72574 133378
rect 71954 133058 71986 133294
rect 72222 133058 72306 133294
rect 72542 133058 72574 133294
rect 71954 73614 72574 133058
rect 71954 73378 71986 73614
rect 72222 73378 72306 73614
rect 72542 73378 72574 73614
rect 71954 73294 72574 73378
rect 71954 73058 71986 73294
rect 72222 73058 72306 73294
rect 72542 73058 72574 73294
rect 71954 13614 72574 73058
rect 71954 13378 71986 13614
rect 72222 13378 72306 13614
rect 72542 13378 72574 13614
rect 71954 13294 72574 13378
rect 71954 13058 71986 13294
rect 72222 13058 72306 13294
rect 72542 13058 72574 13294
rect 41954 -7302 41986 -7066
rect 42222 -7302 42306 -7066
rect 42542 -7302 42574 -7066
rect 41954 -7386 42574 -7302
rect 41954 -7622 41986 -7386
rect 42222 -7622 42306 -7386
rect 42542 -7622 42574 -7386
rect 41954 -7654 42574 -7622
rect 71954 -6106 72574 13058
rect 90794 705798 91414 705830
rect 90794 705562 90826 705798
rect 91062 705562 91146 705798
rect 91382 705562 91414 705798
rect 90794 705478 91414 705562
rect 90794 705242 90826 705478
rect 91062 705242 91146 705478
rect 91382 705242 91414 705478
rect 90794 692454 91414 705242
rect 90794 692218 90826 692454
rect 91062 692218 91146 692454
rect 91382 692218 91414 692454
rect 90794 692134 91414 692218
rect 90794 691898 90826 692134
rect 91062 691898 91146 692134
rect 91382 691898 91414 692134
rect 90794 632454 91414 691898
rect 90794 632218 90826 632454
rect 91062 632218 91146 632454
rect 91382 632218 91414 632454
rect 90794 632134 91414 632218
rect 90794 631898 90826 632134
rect 91062 631898 91146 632134
rect 91382 631898 91414 632134
rect 90794 572454 91414 631898
rect 90794 572218 90826 572454
rect 91062 572218 91146 572454
rect 91382 572218 91414 572454
rect 90794 572134 91414 572218
rect 90794 571898 90826 572134
rect 91062 571898 91146 572134
rect 91382 571898 91414 572134
rect 90794 512454 91414 571898
rect 90794 512218 90826 512454
rect 91062 512218 91146 512454
rect 91382 512218 91414 512454
rect 90794 512134 91414 512218
rect 90794 511898 90826 512134
rect 91062 511898 91146 512134
rect 91382 511898 91414 512134
rect 90794 452454 91414 511898
rect 90794 452218 90826 452454
rect 91062 452218 91146 452454
rect 91382 452218 91414 452454
rect 90794 452134 91414 452218
rect 90794 451898 90826 452134
rect 91062 451898 91146 452134
rect 91382 451898 91414 452134
rect 90794 392454 91414 451898
rect 90794 392218 90826 392454
rect 91062 392218 91146 392454
rect 91382 392218 91414 392454
rect 90794 392134 91414 392218
rect 90794 391898 90826 392134
rect 91062 391898 91146 392134
rect 91382 391898 91414 392134
rect 90794 332454 91414 391898
rect 90794 332218 90826 332454
rect 91062 332218 91146 332454
rect 91382 332218 91414 332454
rect 90794 332134 91414 332218
rect 90794 331898 90826 332134
rect 91062 331898 91146 332134
rect 91382 331898 91414 332134
rect 90794 272454 91414 331898
rect 90794 272218 90826 272454
rect 91062 272218 91146 272454
rect 91382 272218 91414 272454
rect 90794 272134 91414 272218
rect 90794 271898 90826 272134
rect 91062 271898 91146 272134
rect 91382 271898 91414 272134
rect 90794 212454 91414 271898
rect 90794 212218 90826 212454
rect 91062 212218 91146 212454
rect 91382 212218 91414 212454
rect 90794 212134 91414 212218
rect 90794 211898 90826 212134
rect 91062 211898 91146 212134
rect 91382 211898 91414 212134
rect 90794 152454 91414 211898
rect 90794 152218 90826 152454
rect 91062 152218 91146 152454
rect 91382 152218 91414 152454
rect 90794 152134 91414 152218
rect 90794 151898 90826 152134
rect 91062 151898 91146 152134
rect 91382 151898 91414 152134
rect 90794 92454 91414 151898
rect 90794 92218 90826 92454
rect 91062 92218 91146 92454
rect 91382 92218 91414 92454
rect 90794 92134 91414 92218
rect 90794 91898 90826 92134
rect 91062 91898 91146 92134
rect 91382 91898 91414 92134
rect 90794 32454 91414 91898
rect 90794 32218 90826 32454
rect 91062 32218 91146 32454
rect 91382 32218 91414 32454
rect 90794 32134 91414 32218
rect 90794 31898 90826 32134
rect 91062 31898 91146 32134
rect 91382 31898 91414 32134
rect 90794 -1306 91414 31898
rect 90794 -1542 90826 -1306
rect 91062 -1542 91146 -1306
rect 91382 -1542 91414 -1306
rect 90794 -1626 91414 -1542
rect 90794 -1862 90826 -1626
rect 91062 -1862 91146 -1626
rect 91382 -1862 91414 -1626
rect 90794 -1894 91414 -1862
rect 94514 696174 95134 707162
rect 94514 695938 94546 696174
rect 94782 695938 94866 696174
rect 95102 695938 95134 696174
rect 94514 695854 95134 695938
rect 94514 695618 94546 695854
rect 94782 695618 94866 695854
rect 95102 695618 95134 695854
rect 94514 636174 95134 695618
rect 94514 635938 94546 636174
rect 94782 635938 94866 636174
rect 95102 635938 95134 636174
rect 94514 635854 95134 635938
rect 94514 635618 94546 635854
rect 94782 635618 94866 635854
rect 95102 635618 95134 635854
rect 94514 576174 95134 635618
rect 94514 575938 94546 576174
rect 94782 575938 94866 576174
rect 95102 575938 95134 576174
rect 94514 575854 95134 575938
rect 94514 575618 94546 575854
rect 94782 575618 94866 575854
rect 95102 575618 95134 575854
rect 94514 516174 95134 575618
rect 94514 515938 94546 516174
rect 94782 515938 94866 516174
rect 95102 515938 95134 516174
rect 94514 515854 95134 515938
rect 94514 515618 94546 515854
rect 94782 515618 94866 515854
rect 95102 515618 95134 515854
rect 94514 456174 95134 515618
rect 94514 455938 94546 456174
rect 94782 455938 94866 456174
rect 95102 455938 95134 456174
rect 94514 455854 95134 455938
rect 94514 455618 94546 455854
rect 94782 455618 94866 455854
rect 95102 455618 95134 455854
rect 94514 396174 95134 455618
rect 94514 395938 94546 396174
rect 94782 395938 94866 396174
rect 95102 395938 95134 396174
rect 94514 395854 95134 395938
rect 94514 395618 94546 395854
rect 94782 395618 94866 395854
rect 95102 395618 95134 395854
rect 94514 336174 95134 395618
rect 94514 335938 94546 336174
rect 94782 335938 94866 336174
rect 95102 335938 95134 336174
rect 94514 335854 95134 335938
rect 94514 335618 94546 335854
rect 94782 335618 94866 335854
rect 95102 335618 95134 335854
rect 94514 276174 95134 335618
rect 94514 275938 94546 276174
rect 94782 275938 94866 276174
rect 95102 275938 95134 276174
rect 94514 275854 95134 275938
rect 94514 275618 94546 275854
rect 94782 275618 94866 275854
rect 95102 275618 95134 275854
rect 94514 216174 95134 275618
rect 94514 215938 94546 216174
rect 94782 215938 94866 216174
rect 95102 215938 95134 216174
rect 94514 215854 95134 215938
rect 94514 215618 94546 215854
rect 94782 215618 94866 215854
rect 95102 215618 95134 215854
rect 94514 156174 95134 215618
rect 94514 155938 94546 156174
rect 94782 155938 94866 156174
rect 95102 155938 95134 156174
rect 94514 155854 95134 155938
rect 94514 155618 94546 155854
rect 94782 155618 94866 155854
rect 95102 155618 95134 155854
rect 94514 96174 95134 155618
rect 94514 95938 94546 96174
rect 94782 95938 94866 96174
rect 95102 95938 95134 96174
rect 94514 95854 95134 95938
rect 94514 95618 94546 95854
rect 94782 95618 94866 95854
rect 95102 95618 95134 95854
rect 94514 36174 95134 95618
rect 94514 35938 94546 36174
rect 94782 35938 94866 36174
rect 95102 35938 95134 36174
rect 94514 35854 95134 35938
rect 94514 35618 94546 35854
rect 94782 35618 94866 35854
rect 95102 35618 95134 35854
rect 94514 -3226 95134 35618
rect 94514 -3462 94546 -3226
rect 94782 -3462 94866 -3226
rect 95102 -3462 95134 -3226
rect 94514 -3546 95134 -3462
rect 94514 -3782 94546 -3546
rect 94782 -3782 94866 -3546
rect 95102 -3782 95134 -3546
rect 94514 -3814 95134 -3782
rect 98234 699894 98854 709082
rect 98234 699658 98266 699894
rect 98502 699658 98586 699894
rect 98822 699658 98854 699894
rect 98234 699574 98854 699658
rect 98234 699338 98266 699574
rect 98502 699338 98586 699574
rect 98822 699338 98854 699574
rect 98234 639894 98854 699338
rect 98234 639658 98266 639894
rect 98502 639658 98586 639894
rect 98822 639658 98854 639894
rect 98234 639574 98854 639658
rect 98234 639338 98266 639574
rect 98502 639338 98586 639574
rect 98822 639338 98854 639574
rect 98234 579894 98854 639338
rect 98234 579658 98266 579894
rect 98502 579658 98586 579894
rect 98822 579658 98854 579894
rect 98234 579574 98854 579658
rect 98234 579338 98266 579574
rect 98502 579338 98586 579574
rect 98822 579338 98854 579574
rect 98234 519894 98854 579338
rect 98234 519658 98266 519894
rect 98502 519658 98586 519894
rect 98822 519658 98854 519894
rect 98234 519574 98854 519658
rect 98234 519338 98266 519574
rect 98502 519338 98586 519574
rect 98822 519338 98854 519574
rect 98234 459894 98854 519338
rect 98234 459658 98266 459894
rect 98502 459658 98586 459894
rect 98822 459658 98854 459894
rect 98234 459574 98854 459658
rect 98234 459338 98266 459574
rect 98502 459338 98586 459574
rect 98822 459338 98854 459574
rect 98234 399894 98854 459338
rect 98234 399658 98266 399894
rect 98502 399658 98586 399894
rect 98822 399658 98854 399894
rect 98234 399574 98854 399658
rect 98234 399338 98266 399574
rect 98502 399338 98586 399574
rect 98822 399338 98854 399574
rect 98234 339894 98854 399338
rect 98234 339658 98266 339894
rect 98502 339658 98586 339894
rect 98822 339658 98854 339894
rect 98234 339574 98854 339658
rect 98234 339338 98266 339574
rect 98502 339338 98586 339574
rect 98822 339338 98854 339574
rect 98234 279894 98854 339338
rect 98234 279658 98266 279894
rect 98502 279658 98586 279894
rect 98822 279658 98854 279894
rect 98234 279574 98854 279658
rect 98234 279338 98266 279574
rect 98502 279338 98586 279574
rect 98822 279338 98854 279574
rect 98234 219894 98854 279338
rect 98234 219658 98266 219894
rect 98502 219658 98586 219894
rect 98822 219658 98854 219894
rect 98234 219574 98854 219658
rect 98234 219338 98266 219574
rect 98502 219338 98586 219574
rect 98822 219338 98854 219574
rect 98234 159894 98854 219338
rect 98234 159658 98266 159894
rect 98502 159658 98586 159894
rect 98822 159658 98854 159894
rect 98234 159574 98854 159658
rect 98234 159338 98266 159574
rect 98502 159338 98586 159574
rect 98822 159338 98854 159574
rect 98234 99894 98854 159338
rect 98234 99658 98266 99894
rect 98502 99658 98586 99894
rect 98822 99658 98854 99894
rect 98234 99574 98854 99658
rect 98234 99338 98266 99574
rect 98502 99338 98586 99574
rect 98822 99338 98854 99574
rect 98234 39894 98854 99338
rect 98234 39658 98266 39894
rect 98502 39658 98586 39894
rect 98822 39658 98854 39894
rect 98234 39574 98854 39658
rect 98234 39338 98266 39574
rect 98502 39338 98586 39574
rect 98822 39338 98854 39574
rect 98234 -5146 98854 39338
rect 98234 -5382 98266 -5146
rect 98502 -5382 98586 -5146
rect 98822 -5382 98854 -5146
rect 98234 -5466 98854 -5382
rect 98234 -5702 98266 -5466
rect 98502 -5702 98586 -5466
rect 98822 -5702 98854 -5466
rect 98234 -5734 98854 -5702
rect 101954 643614 102574 711002
rect 131954 710598 132574 711590
rect 131954 710362 131986 710598
rect 132222 710362 132306 710598
rect 132542 710362 132574 710598
rect 131954 710278 132574 710362
rect 131954 710042 131986 710278
rect 132222 710042 132306 710278
rect 132542 710042 132574 710278
rect 128234 708678 128854 709670
rect 128234 708442 128266 708678
rect 128502 708442 128586 708678
rect 128822 708442 128854 708678
rect 128234 708358 128854 708442
rect 128234 708122 128266 708358
rect 128502 708122 128586 708358
rect 128822 708122 128854 708358
rect 124514 706758 125134 707750
rect 124514 706522 124546 706758
rect 124782 706522 124866 706758
rect 125102 706522 125134 706758
rect 124514 706438 125134 706522
rect 124514 706202 124546 706438
rect 124782 706202 124866 706438
rect 125102 706202 125134 706438
rect 101954 643378 101986 643614
rect 102222 643378 102306 643614
rect 102542 643378 102574 643614
rect 101954 643294 102574 643378
rect 101954 643058 101986 643294
rect 102222 643058 102306 643294
rect 102542 643058 102574 643294
rect 101954 583614 102574 643058
rect 101954 583378 101986 583614
rect 102222 583378 102306 583614
rect 102542 583378 102574 583614
rect 101954 583294 102574 583378
rect 101954 583058 101986 583294
rect 102222 583058 102306 583294
rect 102542 583058 102574 583294
rect 101954 523614 102574 583058
rect 101954 523378 101986 523614
rect 102222 523378 102306 523614
rect 102542 523378 102574 523614
rect 101954 523294 102574 523378
rect 101954 523058 101986 523294
rect 102222 523058 102306 523294
rect 102542 523058 102574 523294
rect 101954 463614 102574 523058
rect 101954 463378 101986 463614
rect 102222 463378 102306 463614
rect 102542 463378 102574 463614
rect 101954 463294 102574 463378
rect 101954 463058 101986 463294
rect 102222 463058 102306 463294
rect 102542 463058 102574 463294
rect 101954 403614 102574 463058
rect 101954 403378 101986 403614
rect 102222 403378 102306 403614
rect 102542 403378 102574 403614
rect 101954 403294 102574 403378
rect 101954 403058 101986 403294
rect 102222 403058 102306 403294
rect 102542 403058 102574 403294
rect 101954 343614 102574 403058
rect 101954 343378 101986 343614
rect 102222 343378 102306 343614
rect 102542 343378 102574 343614
rect 101954 343294 102574 343378
rect 101954 343058 101986 343294
rect 102222 343058 102306 343294
rect 102542 343058 102574 343294
rect 101954 283614 102574 343058
rect 101954 283378 101986 283614
rect 102222 283378 102306 283614
rect 102542 283378 102574 283614
rect 101954 283294 102574 283378
rect 101954 283058 101986 283294
rect 102222 283058 102306 283294
rect 102542 283058 102574 283294
rect 101954 223614 102574 283058
rect 101954 223378 101986 223614
rect 102222 223378 102306 223614
rect 102542 223378 102574 223614
rect 101954 223294 102574 223378
rect 101954 223058 101986 223294
rect 102222 223058 102306 223294
rect 102542 223058 102574 223294
rect 101954 163614 102574 223058
rect 101954 163378 101986 163614
rect 102222 163378 102306 163614
rect 102542 163378 102574 163614
rect 101954 163294 102574 163378
rect 101954 163058 101986 163294
rect 102222 163058 102306 163294
rect 102542 163058 102574 163294
rect 101954 103614 102574 163058
rect 101954 103378 101986 103614
rect 102222 103378 102306 103614
rect 102542 103378 102574 103614
rect 101954 103294 102574 103378
rect 101954 103058 101986 103294
rect 102222 103058 102306 103294
rect 102542 103058 102574 103294
rect 101954 43614 102574 103058
rect 101954 43378 101986 43614
rect 102222 43378 102306 43614
rect 102542 43378 102574 43614
rect 101954 43294 102574 43378
rect 101954 43058 101986 43294
rect 102222 43058 102306 43294
rect 102542 43058 102574 43294
rect 71954 -6342 71986 -6106
rect 72222 -6342 72306 -6106
rect 72542 -6342 72574 -6106
rect 71954 -6426 72574 -6342
rect 71954 -6662 71986 -6426
rect 72222 -6662 72306 -6426
rect 72542 -6662 72574 -6426
rect 71954 -7654 72574 -6662
rect 101954 -7066 102574 43058
rect 120794 704838 121414 705830
rect 120794 704602 120826 704838
rect 121062 704602 121146 704838
rect 121382 704602 121414 704838
rect 120794 704518 121414 704602
rect 120794 704282 120826 704518
rect 121062 704282 121146 704518
rect 121382 704282 121414 704518
rect 120794 662454 121414 704282
rect 120794 662218 120826 662454
rect 121062 662218 121146 662454
rect 121382 662218 121414 662454
rect 120794 662134 121414 662218
rect 120794 661898 120826 662134
rect 121062 661898 121146 662134
rect 121382 661898 121414 662134
rect 120794 602454 121414 661898
rect 120794 602218 120826 602454
rect 121062 602218 121146 602454
rect 121382 602218 121414 602454
rect 120794 602134 121414 602218
rect 120794 601898 120826 602134
rect 121062 601898 121146 602134
rect 121382 601898 121414 602134
rect 120794 542454 121414 601898
rect 120794 542218 120826 542454
rect 121062 542218 121146 542454
rect 121382 542218 121414 542454
rect 120794 542134 121414 542218
rect 120794 541898 120826 542134
rect 121062 541898 121146 542134
rect 121382 541898 121414 542134
rect 120794 482454 121414 541898
rect 120794 482218 120826 482454
rect 121062 482218 121146 482454
rect 121382 482218 121414 482454
rect 120794 482134 121414 482218
rect 120794 481898 120826 482134
rect 121062 481898 121146 482134
rect 121382 481898 121414 482134
rect 120794 422454 121414 481898
rect 120794 422218 120826 422454
rect 121062 422218 121146 422454
rect 121382 422218 121414 422454
rect 120794 422134 121414 422218
rect 120794 421898 120826 422134
rect 121062 421898 121146 422134
rect 121382 421898 121414 422134
rect 120794 362454 121414 421898
rect 120794 362218 120826 362454
rect 121062 362218 121146 362454
rect 121382 362218 121414 362454
rect 120794 362134 121414 362218
rect 120794 361898 120826 362134
rect 121062 361898 121146 362134
rect 121382 361898 121414 362134
rect 120794 302454 121414 361898
rect 120794 302218 120826 302454
rect 121062 302218 121146 302454
rect 121382 302218 121414 302454
rect 120794 302134 121414 302218
rect 120794 301898 120826 302134
rect 121062 301898 121146 302134
rect 121382 301898 121414 302134
rect 120794 242454 121414 301898
rect 120794 242218 120826 242454
rect 121062 242218 121146 242454
rect 121382 242218 121414 242454
rect 120794 242134 121414 242218
rect 120794 241898 120826 242134
rect 121062 241898 121146 242134
rect 121382 241898 121414 242134
rect 120794 182454 121414 241898
rect 120794 182218 120826 182454
rect 121062 182218 121146 182454
rect 121382 182218 121414 182454
rect 120794 182134 121414 182218
rect 120794 181898 120826 182134
rect 121062 181898 121146 182134
rect 121382 181898 121414 182134
rect 120794 122454 121414 181898
rect 120794 122218 120826 122454
rect 121062 122218 121146 122454
rect 121382 122218 121414 122454
rect 120794 122134 121414 122218
rect 120794 121898 120826 122134
rect 121062 121898 121146 122134
rect 121382 121898 121414 122134
rect 120794 62454 121414 121898
rect 120794 62218 120826 62454
rect 121062 62218 121146 62454
rect 121382 62218 121414 62454
rect 120794 62134 121414 62218
rect 120794 61898 120826 62134
rect 121062 61898 121146 62134
rect 121382 61898 121414 62134
rect 120794 2454 121414 61898
rect 120794 2218 120826 2454
rect 121062 2218 121146 2454
rect 121382 2218 121414 2454
rect 120794 2134 121414 2218
rect 120794 1898 120826 2134
rect 121062 1898 121146 2134
rect 121382 1898 121414 2134
rect 120794 -346 121414 1898
rect 120794 -582 120826 -346
rect 121062 -582 121146 -346
rect 121382 -582 121414 -346
rect 120794 -666 121414 -582
rect 120794 -902 120826 -666
rect 121062 -902 121146 -666
rect 121382 -902 121414 -666
rect 120794 -1894 121414 -902
rect 124514 666174 125134 706202
rect 124514 665938 124546 666174
rect 124782 665938 124866 666174
rect 125102 665938 125134 666174
rect 124514 665854 125134 665938
rect 124514 665618 124546 665854
rect 124782 665618 124866 665854
rect 125102 665618 125134 665854
rect 124514 606174 125134 665618
rect 124514 605938 124546 606174
rect 124782 605938 124866 606174
rect 125102 605938 125134 606174
rect 124514 605854 125134 605938
rect 124514 605618 124546 605854
rect 124782 605618 124866 605854
rect 125102 605618 125134 605854
rect 124514 546174 125134 605618
rect 124514 545938 124546 546174
rect 124782 545938 124866 546174
rect 125102 545938 125134 546174
rect 124514 545854 125134 545938
rect 124514 545618 124546 545854
rect 124782 545618 124866 545854
rect 125102 545618 125134 545854
rect 124514 486174 125134 545618
rect 124514 485938 124546 486174
rect 124782 485938 124866 486174
rect 125102 485938 125134 486174
rect 124514 485854 125134 485938
rect 124514 485618 124546 485854
rect 124782 485618 124866 485854
rect 125102 485618 125134 485854
rect 124514 426174 125134 485618
rect 124514 425938 124546 426174
rect 124782 425938 124866 426174
rect 125102 425938 125134 426174
rect 124514 425854 125134 425938
rect 124514 425618 124546 425854
rect 124782 425618 124866 425854
rect 125102 425618 125134 425854
rect 124514 366174 125134 425618
rect 124514 365938 124546 366174
rect 124782 365938 124866 366174
rect 125102 365938 125134 366174
rect 124514 365854 125134 365938
rect 124514 365618 124546 365854
rect 124782 365618 124866 365854
rect 125102 365618 125134 365854
rect 124514 306174 125134 365618
rect 124514 305938 124546 306174
rect 124782 305938 124866 306174
rect 125102 305938 125134 306174
rect 124514 305854 125134 305938
rect 124514 305618 124546 305854
rect 124782 305618 124866 305854
rect 125102 305618 125134 305854
rect 124514 246174 125134 305618
rect 124514 245938 124546 246174
rect 124782 245938 124866 246174
rect 125102 245938 125134 246174
rect 124514 245854 125134 245938
rect 124514 245618 124546 245854
rect 124782 245618 124866 245854
rect 125102 245618 125134 245854
rect 124514 186174 125134 245618
rect 124514 185938 124546 186174
rect 124782 185938 124866 186174
rect 125102 185938 125134 186174
rect 124514 185854 125134 185938
rect 124514 185618 124546 185854
rect 124782 185618 124866 185854
rect 125102 185618 125134 185854
rect 124514 126174 125134 185618
rect 124514 125938 124546 126174
rect 124782 125938 124866 126174
rect 125102 125938 125134 126174
rect 124514 125854 125134 125938
rect 124514 125618 124546 125854
rect 124782 125618 124866 125854
rect 125102 125618 125134 125854
rect 124514 66174 125134 125618
rect 124514 65938 124546 66174
rect 124782 65938 124866 66174
rect 125102 65938 125134 66174
rect 124514 65854 125134 65938
rect 124514 65618 124546 65854
rect 124782 65618 124866 65854
rect 125102 65618 125134 65854
rect 124514 6174 125134 65618
rect 124514 5938 124546 6174
rect 124782 5938 124866 6174
rect 125102 5938 125134 6174
rect 124514 5854 125134 5938
rect 124514 5618 124546 5854
rect 124782 5618 124866 5854
rect 125102 5618 125134 5854
rect 124514 -2266 125134 5618
rect 124514 -2502 124546 -2266
rect 124782 -2502 124866 -2266
rect 125102 -2502 125134 -2266
rect 124514 -2586 125134 -2502
rect 124514 -2822 124546 -2586
rect 124782 -2822 124866 -2586
rect 125102 -2822 125134 -2586
rect 124514 -3814 125134 -2822
rect 128234 669894 128854 708122
rect 128234 669658 128266 669894
rect 128502 669658 128586 669894
rect 128822 669658 128854 669894
rect 128234 669574 128854 669658
rect 128234 669338 128266 669574
rect 128502 669338 128586 669574
rect 128822 669338 128854 669574
rect 128234 609894 128854 669338
rect 128234 609658 128266 609894
rect 128502 609658 128586 609894
rect 128822 609658 128854 609894
rect 128234 609574 128854 609658
rect 128234 609338 128266 609574
rect 128502 609338 128586 609574
rect 128822 609338 128854 609574
rect 128234 549894 128854 609338
rect 128234 549658 128266 549894
rect 128502 549658 128586 549894
rect 128822 549658 128854 549894
rect 128234 549574 128854 549658
rect 128234 549338 128266 549574
rect 128502 549338 128586 549574
rect 128822 549338 128854 549574
rect 128234 489894 128854 549338
rect 128234 489658 128266 489894
rect 128502 489658 128586 489894
rect 128822 489658 128854 489894
rect 128234 489574 128854 489658
rect 128234 489338 128266 489574
rect 128502 489338 128586 489574
rect 128822 489338 128854 489574
rect 128234 429894 128854 489338
rect 128234 429658 128266 429894
rect 128502 429658 128586 429894
rect 128822 429658 128854 429894
rect 128234 429574 128854 429658
rect 128234 429338 128266 429574
rect 128502 429338 128586 429574
rect 128822 429338 128854 429574
rect 128234 369894 128854 429338
rect 128234 369658 128266 369894
rect 128502 369658 128586 369894
rect 128822 369658 128854 369894
rect 128234 369574 128854 369658
rect 128234 369338 128266 369574
rect 128502 369338 128586 369574
rect 128822 369338 128854 369574
rect 128234 309894 128854 369338
rect 128234 309658 128266 309894
rect 128502 309658 128586 309894
rect 128822 309658 128854 309894
rect 128234 309574 128854 309658
rect 128234 309338 128266 309574
rect 128502 309338 128586 309574
rect 128822 309338 128854 309574
rect 128234 249894 128854 309338
rect 128234 249658 128266 249894
rect 128502 249658 128586 249894
rect 128822 249658 128854 249894
rect 128234 249574 128854 249658
rect 128234 249338 128266 249574
rect 128502 249338 128586 249574
rect 128822 249338 128854 249574
rect 128234 189894 128854 249338
rect 128234 189658 128266 189894
rect 128502 189658 128586 189894
rect 128822 189658 128854 189894
rect 128234 189574 128854 189658
rect 128234 189338 128266 189574
rect 128502 189338 128586 189574
rect 128822 189338 128854 189574
rect 128234 129894 128854 189338
rect 128234 129658 128266 129894
rect 128502 129658 128586 129894
rect 128822 129658 128854 129894
rect 128234 129574 128854 129658
rect 128234 129338 128266 129574
rect 128502 129338 128586 129574
rect 128822 129338 128854 129574
rect 128234 69894 128854 129338
rect 128234 69658 128266 69894
rect 128502 69658 128586 69894
rect 128822 69658 128854 69894
rect 128234 69574 128854 69658
rect 128234 69338 128266 69574
rect 128502 69338 128586 69574
rect 128822 69338 128854 69574
rect 128234 9894 128854 69338
rect 128234 9658 128266 9894
rect 128502 9658 128586 9894
rect 128822 9658 128854 9894
rect 128234 9574 128854 9658
rect 128234 9338 128266 9574
rect 128502 9338 128586 9574
rect 128822 9338 128854 9574
rect 128234 -4186 128854 9338
rect 128234 -4422 128266 -4186
rect 128502 -4422 128586 -4186
rect 128822 -4422 128854 -4186
rect 128234 -4506 128854 -4422
rect 128234 -4742 128266 -4506
rect 128502 -4742 128586 -4506
rect 128822 -4742 128854 -4506
rect 128234 -5734 128854 -4742
rect 131954 673614 132574 710042
rect 161954 711558 162574 711590
rect 161954 711322 161986 711558
rect 162222 711322 162306 711558
rect 162542 711322 162574 711558
rect 161954 711238 162574 711322
rect 161954 711002 161986 711238
rect 162222 711002 162306 711238
rect 162542 711002 162574 711238
rect 158234 709638 158854 709670
rect 158234 709402 158266 709638
rect 158502 709402 158586 709638
rect 158822 709402 158854 709638
rect 158234 709318 158854 709402
rect 158234 709082 158266 709318
rect 158502 709082 158586 709318
rect 158822 709082 158854 709318
rect 154514 707718 155134 707750
rect 154514 707482 154546 707718
rect 154782 707482 154866 707718
rect 155102 707482 155134 707718
rect 154514 707398 155134 707482
rect 154514 707162 154546 707398
rect 154782 707162 154866 707398
rect 155102 707162 155134 707398
rect 131954 673378 131986 673614
rect 132222 673378 132306 673614
rect 132542 673378 132574 673614
rect 131954 673294 132574 673378
rect 131954 673058 131986 673294
rect 132222 673058 132306 673294
rect 132542 673058 132574 673294
rect 131954 613614 132574 673058
rect 131954 613378 131986 613614
rect 132222 613378 132306 613614
rect 132542 613378 132574 613614
rect 131954 613294 132574 613378
rect 131954 613058 131986 613294
rect 132222 613058 132306 613294
rect 132542 613058 132574 613294
rect 131954 553614 132574 613058
rect 131954 553378 131986 553614
rect 132222 553378 132306 553614
rect 132542 553378 132574 553614
rect 131954 553294 132574 553378
rect 131954 553058 131986 553294
rect 132222 553058 132306 553294
rect 132542 553058 132574 553294
rect 131954 493614 132574 553058
rect 131954 493378 131986 493614
rect 132222 493378 132306 493614
rect 132542 493378 132574 493614
rect 131954 493294 132574 493378
rect 131954 493058 131986 493294
rect 132222 493058 132306 493294
rect 132542 493058 132574 493294
rect 131954 433614 132574 493058
rect 131954 433378 131986 433614
rect 132222 433378 132306 433614
rect 132542 433378 132574 433614
rect 131954 433294 132574 433378
rect 131954 433058 131986 433294
rect 132222 433058 132306 433294
rect 132542 433058 132574 433294
rect 131954 373614 132574 433058
rect 131954 373378 131986 373614
rect 132222 373378 132306 373614
rect 132542 373378 132574 373614
rect 131954 373294 132574 373378
rect 131954 373058 131986 373294
rect 132222 373058 132306 373294
rect 132542 373058 132574 373294
rect 131954 313614 132574 373058
rect 131954 313378 131986 313614
rect 132222 313378 132306 313614
rect 132542 313378 132574 313614
rect 131954 313294 132574 313378
rect 131954 313058 131986 313294
rect 132222 313058 132306 313294
rect 132542 313058 132574 313294
rect 131954 253614 132574 313058
rect 131954 253378 131986 253614
rect 132222 253378 132306 253614
rect 132542 253378 132574 253614
rect 131954 253294 132574 253378
rect 131954 253058 131986 253294
rect 132222 253058 132306 253294
rect 132542 253058 132574 253294
rect 131954 193614 132574 253058
rect 131954 193378 131986 193614
rect 132222 193378 132306 193614
rect 132542 193378 132574 193614
rect 131954 193294 132574 193378
rect 131954 193058 131986 193294
rect 132222 193058 132306 193294
rect 132542 193058 132574 193294
rect 131954 133614 132574 193058
rect 131954 133378 131986 133614
rect 132222 133378 132306 133614
rect 132542 133378 132574 133614
rect 131954 133294 132574 133378
rect 131954 133058 131986 133294
rect 132222 133058 132306 133294
rect 132542 133058 132574 133294
rect 131954 73614 132574 133058
rect 131954 73378 131986 73614
rect 132222 73378 132306 73614
rect 132542 73378 132574 73614
rect 131954 73294 132574 73378
rect 131954 73058 131986 73294
rect 132222 73058 132306 73294
rect 132542 73058 132574 73294
rect 131954 13614 132574 73058
rect 131954 13378 131986 13614
rect 132222 13378 132306 13614
rect 132542 13378 132574 13614
rect 131954 13294 132574 13378
rect 131954 13058 131986 13294
rect 132222 13058 132306 13294
rect 132542 13058 132574 13294
rect 101954 -7302 101986 -7066
rect 102222 -7302 102306 -7066
rect 102542 -7302 102574 -7066
rect 101954 -7386 102574 -7302
rect 101954 -7622 101986 -7386
rect 102222 -7622 102306 -7386
rect 102542 -7622 102574 -7386
rect 101954 -7654 102574 -7622
rect 131954 -6106 132574 13058
rect 150794 705798 151414 705830
rect 150794 705562 150826 705798
rect 151062 705562 151146 705798
rect 151382 705562 151414 705798
rect 150794 705478 151414 705562
rect 150794 705242 150826 705478
rect 151062 705242 151146 705478
rect 151382 705242 151414 705478
rect 150794 692454 151414 705242
rect 150794 692218 150826 692454
rect 151062 692218 151146 692454
rect 151382 692218 151414 692454
rect 150794 692134 151414 692218
rect 150794 691898 150826 692134
rect 151062 691898 151146 692134
rect 151382 691898 151414 692134
rect 150794 632454 151414 691898
rect 150794 632218 150826 632454
rect 151062 632218 151146 632454
rect 151382 632218 151414 632454
rect 150794 632134 151414 632218
rect 150794 631898 150826 632134
rect 151062 631898 151146 632134
rect 151382 631898 151414 632134
rect 150794 572454 151414 631898
rect 150794 572218 150826 572454
rect 151062 572218 151146 572454
rect 151382 572218 151414 572454
rect 150794 572134 151414 572218
rect 150794 571898 150826 572134
rect 151062 571898 151146 572134
rect 151382 571898 151414 572134
rect 150794 512454 151414 571898
rect 150794 512218 150826 512454
rect 151062 512218 151146 512454
rect 151382 512218 151414 512454
rect 150794 512134 151414 512218
rect 150794 511898 150826 512134
rect 151062 511898 151146 512134
rect 151382 511898 151414 512134
rect 150794 452454 151414 511898
rect 150794 452218 150826 452454
rect 151062 452218 151146 452454
rect 151382 452218 151414 452454
rect 150794 452134 151414 452218
rect 150794 451898 150826 452134
rect 151062 451898 151146 452134
rect 151382 451898 151414 452134
rect 150794 392454 151414 451898
rect 150794 392218 150826 392454
rect 151062 392218 151146 392454
rect 151382 392218 151414 392454
rect 150794 392134 151414 392218
rect 150794 391898 150826 392134
rect 151062 391898 151146 392134
rect 151382 391898 151414 392134
rect 150794 332454 151414 391898
rect 150794 332218 150826 332454
rect 151062 332218 151146 332454
rect 151382 332218 151414 332454
rect 150794 332134 151414 332218
rect 150794 331898 150826 332134
rect 151062 331898 151146 332134
rect 151382 331898 151414 332134
rect 150794 272454 151414 331898
rect 150794 272218 150826 272454
rect 151062 272218 151146 272454
rect 151382 272218 151414 272454
rect 150794 272134 151414 272218
rect 150794 271898 150826 272134
rect 151062 271898 151146 272134
rect 151382 271898 151414 272134
rect 150794 212454 151414 271898
rect 150794 212218 150826 212454
rect 151062 212218 151146 212454
rect 151382 212218 151414 212454
rect 150794 212134 151414 212218
rect 150794 211898 150826 212134
rect 151062 211898 151146 212134
rect 151382 211898 151414 212134
rect 150794 152454 151414 211898
rect 150794 152218 150826 152454
rect 151062 152218 151146 152454
rect 151382 152218 151414 152454
rect 150794 152134 151414 152218
rect 150794 151898 150826 152134
rect 151062 151898 151146 152134
rect 151382 151898 151414 152134
rect 150794 92454 151414 151898
rect 150794 92218 150826 92454
rect 151062 92218 151146 92454
rect 151382 92218 151414 92454
rect 150794 92134 151414 92218
rect 150794 91898 150826 92134
rect 151062 91898 151146 92134
rect 151382 91898 151414 92134
rect 150794 32454 151414 91898
rect 150794 32218 150826 32454
rect 151062 32218 151146 32454
rect 151382 32218 151414 32454
rect 150794 32134 151414 32218
rect 150794 31898 150826 32134
rect 151062 31898 151146 32134
rect 151382 31898 151414 32134
rect 150794 -1306 151414 31898
rect 150794 -1542 150826 -1306
rect 151062 -1542 151146 -1306
rect 151382 -1542 151414 -1306
rect 150794 -1626 151414 -1542
rect 150794 -1862 150826 -1626
rect 151062 -1862 151146 -1626
rect 151382 -1862 151414 -1626
rect 150794 -1894 151414 -1862
rect 154514 696174 155134 707162
rect 154514 695938 154546 696174
rect 154782 695938 154866 696174
rect 155102 695938 155134 696174
rect 154514 695854 155134 695938
rect 154514 695618 154546 695854
rect 154782 695618 154866 695854
rect 155102 695618 155134 695854
rect 154514 636174 155134 695618
rect 154514 635938 154546 636174
rect 154782 635938 154866 636174
rect 155102 635938 155134 636174
rect 154514 635854 155134 635938
rect 154514 635618 154546 635854
rect 154782 635618 154866 635854
rect 155102 635618 155134 635854
rect 154514 576174 155134 635618
rect 154514 575938 154546 576174
rect 154782 575938 154866 576174
rect 155102 575938 155134 576174
rect 154514 575854 155134 575938
rect 154514 575618 154546 575854
rect 154782 575618 154866 575854
rect 155102 575618 155134 575854
rect 154514 516174 155134 575618
rect 154514 515938 154546 516174
rect 154782 515938 154866 516174
rect 155102 515938 155134 516174
rect 154514 515854 155134 515938
rect 154514 515618 154546 515854
rect 154782 515618 154866 515854
rect 155102 515618 155134 515854
rect 154514 456174 155134 515618
rect 154514 455938 154546 456174
rect 154782 455938 154866 456174
rect 155102 455938 155134 456174
rect 154514 455854 155134 455938
rect 154514 455618 154546 455854
rect 154782 455618 154866 455854
rect 155102 455618 155134 455854
rect 154514 396174 155134 455618
rect 154514 395938 154546 396174
rect 154782 395938 154866 396174
rect 155102 395938 155134 396174
rect 154514 395854 155134 395938
rect 154514 395618 154546 395854
rect 154782 395618 154866 395854
rect 155102 395618 155134 395854
rect 154514 336174 155134 395618
rect 154514 335938 154546 336174
rect 154782 335938 154866 336174
rect 155102 335938 155134 336174
rect 154514 335854 155134 335938
rect 154514 335618 154546 335854
rect 154782 335618 154866 335854
rect 155102 335618 155134 335854
rect 154514 276174 155134 335618
rect 154514 275938 154546 276174
rect 154782 275938 154866 276174
rect 155102 275938 155134 276174
rect 154514 275854 155134 275938
rect 154514 275618 154546 275854
rect 154782 275618 154866 275854
rect 155102 275618 155134 275854
rect 154514 216174 155134 275618
rect 154514 215938 154546 216174
rect 154782 215938 154866 216174
rect 155102 215938 155134 216174
rect 154514 215854 155134 215938
rect 154514 215618 154546 215854
rect 154782 215618 154866 215854
rect 155102 215618 155134 215854
rect 154514 156174 155134 215618
rect 154514 155938 154546 156174
rect 154782 155938 154866 156174
rect 155102 155938 155134 156174
rect 154514 155854 155134 155938
rect 154514 155618 154546 155854
rect 154782 155618 154866 155854
rect 155102 155618 155134 155854
rect 154514 96174 155134 155618
rect 154514 95938 154546 96174
rect 154782 95938 154866 96174
rect 155102 95938 155134 96174
rect 154514 95854 155134 95938
rect 154514 95618 154546 95854
rect 154782 95618 154866 95854
rect 155102 95618 155134 95854
rect 154514 36174 155134 95618
rect 154514 35938 154546 36174
rect 154782 35938 154866 36174
rect 155102 35938 155134 36174
rect 154514 35854 155134 35938
rect 154514 35618 154546 35854
rect 154782 35618 154866 35854
rect 155102 35618 155134 35854
rect 154514 -3226 155134 35618
rect 154514 -3462 154546 -3226
rect 154782 -3462 154866 -3226
rect 155102 -3462 155134 -3226
rect 154514 -3546 155134 -3462
rect 154514 -3782 154546 -3546
rect 154782 -3782 154866 -3546
rect 155102 -3782 155134 -3546
rect 154514 -3814 155134 -3782
rect 158234 699894 158854 709082
rect 158234 699658 158266 699894
rect 158502 699658 158586 699894
rect 158822 699658 158854 699894
rect 158234 699574 158854 699658
rect 158234 699338 158266 699574
rect 158502 699338 158586 699574
rect 158822 699338 158854 699574
rect 158234 639894 158854 699338
rect 158234 639658 158266 639894
rect 158502 639658 158586 639894
rect 158822 639658 158854 639894
rect 158234 639574 158854 639658
rect 158234 639338 158266 639574
rect 158502 639338 158586 639574
rect 158822 639338 158854 639574
rect 158234 579894 158854 639338
rect 158234 579658 158266 579894
rect 158502 579658 158586 579894
rect 158822 579658 158854 579894
rect 158234 579574 158854 579658
rect 158234 579338 158266 579574
rect 158502 579338 158586 579574
rect 158822 579338 158854 579574
rect 158234 519894 158854 579338
rect 158234 519658 158266 519894
rect 158502 519658 158586 519894
rect 158822 519658 158854 519894
rect 158234 519574 158854 519658
rect 158234 519338 158266 519574
rect 158502 519338 158586 519574
rect 158822 519338 158854 519574
rect 158234 459894 158854 519338
rect 158234 459658 158266 459894
rect 158502 459658 158586 459894
rect 158822 459658 158854 459894
rect 158234 459574 158854 459658
rect 158234 459338 158266 459574
rect 158502 459338 158586 459574
rect 158822 459338 158854 459574
rect 158234 399894 158854 459338
rect 158234 399658 158266 399894
rect 158502 399658 158586 399894
rect 158822 399658 158854 399894
rect 158234 399574 158854 399658
rect 158234 399338 158266 399574
rect 158502 399338 158586 399574
rect 158822 399338 158854 399574
rect 158234 339894 158854 399338
rect 158234 339658 158266 339894
rect 158502 339658 158586 339894
rect 158822 339658 158854 339894
rect 158234 339574 158854 339658
rect 158234 339338 158266 339574
rect 158502 339338 158586 339574
rect 158822 339338 158854 339574
rect 158234 279894 158854 339338
rect 158234 279658 158266 279894
rect 158502 279658 158586 279894
rect 158822 279658 158854 279894
rect 158234 279574 158854 279658
rect 158234 279338 158266 279574
rect 158502 279338 158586 279574
rect 158822 279338 158854 279574
rect 158234 219894 158854 279338
rect 158234 219658 158266 219894
rect 158502 219658 158586 219894
rect 158822 219658 158854 219894
rect 158234 219574 158854 219658
rect 158234 219338 158266 219574
rect 158502 219338 158586 219574
rect 158822 219338 158854 219574
rect 158234 159894 158854 219338
rect 158234 159658 158266 159894
rect 158502 159658 158586 159894
rect 158822 159658 158854 159894
rect 158234 159574 158854 159658
rect 158234 159338 158266 159574
rect 158502 159338 158586 159574
rect 158822 159338 158854 159574
rect 158234 99894 158854 159338
rect 158234 99658 158266 99894
rect 158502 99658 158586 99894
rect 158822 99658 158854 99894
rect 158234 99574 158854 99658
rect 158234 99338 158266 99574
rect 158502 99338 158586 99574
rect 158822 99338 158854 99574
rect 158234 39894 158854 99338
rect 158234 39658 158266 39894
rect 158502 39658 158586 39894
rect 158822 39658 158854 39894
rect 158234 39574 158854 39658
rect 158234 39338 158266 39574
rect 158502 39338 158586 39574
rect 158822 39338 158854 39574
rect 158234 -5146 158854 39338
rect 158234 -5382 158266 -5146
rect 158502 -5382 158586 -5146
rect 158822 -5382 158854 -5146
rect 158234 -5466 158854 -5382
rect 158234 -5702 158266 -5466
rect 158502 -5702 158586 -5466
rect 158822 -5702 158854 -5466
rect 158234 -5734 158854 -5702
rect 161954 643614 162574 711002
rect 191954 710598 192574 711590
rect 191954 710362 191986 710598
rect 192222 710362 192306 710598
rect 192542 710362 192574 710598
rect 191954 710278 192574 710362
rect 191954 710042 191986 710278
rect 192222 710042 192306 710278
rect 192542 710042 192574 710278
rect 188234 708678 188854 709670
rect 188234 708442 188266 708678
rect 188502 708442 188586 708678
rect 188822 708442 188854 708678
rect 188234 708358 188854 708442
rect 188234 708122 188266 708358
rect 188502 708122 188586 708358
rect 188822 708122 188854 708358
rect 184514 706758 185134 707750
rect 184514 706522 184546 706758
rect 184782 706522 184866 706758
rect 185102 706522 185134 706758
rect 184514 706438 185134 706522
rect 184514 706202 184546 706438
rect 184782 706202 184866 706438
rect 185102 706202 185134 706438
rect 161954 643378 161986 643614
rect 162222 643378 162306 643614
rect 162542 643378 162574 643614
rect 161954 643294 162574 643378
rect 161954 643058 161986 643294
rect 162222 643058 162306 643294
rect 162542 643058 162574 643294
rect 161954 583614 162574 643058
rect 161954 583378 161986 583614
rect 162222 583378 162306 583614
rect 162542 583378 162574 583614
rect 161954 583294 162574 583378
rect 161954 583058 161986 583294
rect 162222 583058 162306 583294
rect 162542 583058 162574 583294
rect 161954 523614 162574 583058
rect 161954 523378 161986 523614
rect 162222 523378 162306 523614
rect 162542 523378 162574 523614
rect 161954 523294 162574 523378
rect 161954 523058 161986 523294
rect 162222 523058 162306 523294
rect 162542 523058 162574 523294
rect 161954 463614 162574 523058
rect 161954 463378 161986 463614
rect 162222 463378 162306 463614
rect 162542 463378 162574 463614
rect 161954 463294 162574 463378
rect 161954 463058 161986 463294
rect 162222 463058 162306 463294
rect 162542 463058 162574 463294
rect 161954 403614 162574 463058
rect 161954 403378 161986 403614
rect 162222 403378 162306 403614
rect 162542 403378 162574 403614
rect 161954 403294 162574 403378
rect 161954 403058 161986 403294
rect 162222 403058 162306 403294
rect 162542 403058 162574 403294
rect 161954 343614 162574 403058
rect 161954 343378 161986 343614
rect 162222 343378 162306 343614
rect 162542 343378 162574 343614
rect 161954 343294 162574 343378
rect 161954 343058 161986 343294
rect 162222 343058 162306 343294
rect 162542 343058 162574 343294
rect 161954 283614 162574 343058
rect 161954 283378 161986 283614
rect 162222 283378 162306 283614
rect 162542 283378 162574 283614
rect 161954 283294 162574 283378
rect 161954 283058 161986 283294
rect 162222 283058 162306 283294
rect 162542 283058 162574 283294
rect 161954 223614 162574 283058
rect 161954 223378 161986 223614
rect 162222 223378 162306 223614
rect 162542 223378 162574 223614
rect 161954 223294 162574 223378
rect 161954 223058 161986 223294
rect 162222 223058 162306 223294
rect 162542 223058 162574 223294
rect 161954 163614 162574 223058
rect 161954 163378 161986 163614
rect 162222 163378 162306 163614
rect 162542 163378 162574 163614
rect 161954 163294 162574 163378
rect 161954 163058 161986 163294
rect 162222 163058 162306 163294
rect 162542 163058 162574 163294
rect 161954 103614 162574 163058
rect 161954 103378 161986 103614
rect 162222 103378 162306 103614
rect 162542 103378 162574 103614
rect 161954 103294 162574 103378
rect 161954 103058 161986 103294
rect 162222 103058 162306 103294
rect 162542 103058 162574 103294
rect 161954 43614 162574 103058
rect 161954 43378 161986 43614
rect 162222 43378 162306 43614
rect 162542 43378 162574 43614
rect 161954 43294 162574 43378
rect 161954 43058 161986 43294
rect 162222 43058 162306 43294
rect 162542 43058 162574 43294
rect 131954 -6342 131986 -6106
rect 132222 -6342 132306 -6106
rect 132542 -6342 132574 -6106
rect 131954 -6426 132574 -6342
rect 131954 -6662 131986 -6426
rect 132222 -6662 132306 -6426
rect 132542 -6662 132574 -6426
rect 131954 -7654 132574 -6662
rect 161954 -7066 162574 43058
rect 180794 704838 181414 705830
rect 180794 704602 180826 704838
rect 181062 704602 181146 704838
rect 181382 704602 181414 704838
rect 180794 704518 181414 704602
rect 180794 704282 180826 704518
rect 181062 704282 181146 704518
rect 181382 704282 181414 704518
rect 180794 662454 181414 704282
rect 180794 662218 180826 662454
rect 181062 662218 181146 662454
rect 181382 662218 181414 662454
rect 180794 662134 181414 662218
rect 180794 661898 180826 662134
rect 181062 661898 181146 662134
rect 181382 661898 181414 662134
rect 180794 602454 181414 661898
rect 180794 602218 180826 602454
rect 181062 602218 181146 602454
rect 181382 602218 181414 602454
rect 180794 602134 181414 602218
rect 180794 601898 180826 602134
rect 181062 601898 181146 602134
rect 181382 601898 181414 602134
rect 180794 542454 181414 601898
rect 180794 542218 180826 542454
rect 181062 542218 181146 542454
rect 181382 542218 181414 542454
rect 180794 542134 181414 542218
rect 180794 541898 180826 542134
rect 181062 541898 181146 542134
rect 181382 541898 181414 542134
rect 180794 482454 181414 541898
rect 180794 482218 180826 482454
rect 181062 482218 181146 482454
rect 181382 482218 181414 482454
rect 180794 482134 181414 482218
rect 180794 481898 180826 482134
rect 181062 481898 181146 482134
rect 181382 481898 181414 482134
rect 180794 422454 181414 481898
rect 180794 422218 180826 422454
rect 181062 422218 181146 422454
rect 181382 422218 181414 422454
rect 180794 422134 181414 422218
rect 180794 421898 180826 422134
rect 181062 421898 181146 422134
rect 181382 421898 181414 422134
rect 180794 362454 181414 421898
rect 180794 362218 180826 362454
rect 181062 362218 181146 362454
rect 181382 362218 181414 362454
rect 180794 362134 181414 362218
rect 180794 361898 180826 362134
rect 181062 361898 181146 362134
rect 181382 361898 181414 362134
rect 180794 302454 181414 361898
rect 180794 302218 180826 302454
rect 181062 302218 181146 302454
rect 181382 302218 181414 302454
rect 180794 302134 181414 302218
rect 180794 301898 180826 302134
rect 181062 301898 181146 302134
rect 181382 301898 181414 302134
rect 180794 242454 181414 301898
rect 180794 242218 180826 242454
rect 181062 242218 181146 242454
rect 181382 242218 181414 242454
rect 180794 242134 181414 242218
rect 180794 241898 180826 242134
rect 181062 241898 181146 242134
rect 181382 241898 181414 242134
rect 180794 182454 181414 241898
rect 180794 182218 180826 182454
rect 181062 182218 181146 182454
rect 181382 182218 181414 182454
rect 180794 182134 181414 182218
rect 180794 181898 180826 182134
rect 181062 181898 181146 182134
rect 181382 181898 181414 182134
rect 180794 122454 181414 181898
rect 180794 122218 180826 122454
rect 181062 122218 181146 122454
rect 181382 122218 181414 122454
rect 180794 122134 181414 122218
rect 180794 121898 180826 122134
rect 181062 121898 181146 122134
rect 181382 121898 181414 122134
rect 180794 62454 181414 121898
rect 180794 62218 180826 62454
rect 181062 62218 181146 62454
rect 181382 62218 181414 62454
rect 180794 62134 181414 62218
rect 180794 61898 180826 62134
rect 181062 61898 181146 62134
rect 181382 61898 181414 62134
rect 180794 2454 181414 61898
rect 180794 2218 180826 2454
rect 181062 2218 181146 2454
rect 181382 2218 181414 2454
rect 180794 2134 181414 2218
rect 180794 1898 180826 2134
rect 181062 1898 181146 2134
rect 181382 1898 181414 2134
rect 180794 -346 181414 1898
rect 180794 -582 180826 -346
rect 181062 -582 181146 -346
rect 181382 -582 181414 -346
rect 180794 -666 181414 -582
rect 180794 -902 180826 -666
rect 181062 -902 181146 -666
rect 181382 -902 181414 -666
rect 180794 -1894 181414 -902
rect 184514 666174 185134 706202
rect 184514 665938 184546 666174
rect 184782 665938 184866 666174
rect 185102 665938 185134 666174
rect 184514 665854 185134 665938
rect 184514 665618 184546 665854
rect 184782 665618 184866 665854
rect 185102 665618 185134 665854
rect 184514 606174 185134 665618
rect 184514 605938 184546 606174
rect 184782 605938 184866 606174
rect 185102 605938 185134 606174
rect 184514 605854 185134 605938
rect 184514 605618 184546 605854
rect 184782 605618 184866 605854
rect 185102 605618 185134 605854
rect 184514 546174 185134 605618
rect 184514 545938 184546 546174
rect 184782 545938 184866 546174
rect 185102 545938 185134 546174
rect 184514 545854 185134 545938
rect 184514 545618 184546 545854
rect 184782 545618 184866 545854
rect 185102 545618 185134 545854
rect 184514 486174 185134 545618
rect 184514 485938 184546 486174
rect 184782 485938 184866 486174
rect 185102 485938 185134 486174
rect 184514 485854 185134 485938
rect 184514 485618 184546 485854
rect 184782 485618 184866 485854
rect 185102 485618 185134 485854
rect 184514 426174 185134 485618
rect 184514 425938 184546 426174
rect 184782 425938 184866 426174
rect 185102 425938 185134 426174
rect 184514 425854 185134 425938
rect 184514 425618 184546 425854
rect 184782 425618 184866 425854
rect 185102 425618 185134 425854
rect 184514 366174 185134 425618
rect 184514 365938 184546 366174
rect 184782 365938 184866 366174
rect 185102 365938 185134 366174
rect 184514 365854 185134 365938
rect 184514 365618 184546 365854
rect 184782 365618 184866 365854
rect 185102 365618 185134 365854
rect 184514 306174 185134 365618
rect 184514 305938 184546 306174
rect 184782 305938 184866 306174
rect 185102 305938 185134 306174
rect 184514 305854 185134 305938
rect 184514 305618 184546 305854
rect 184782 305618 184866 305854
rect 185102 305618 185134 305854
rect 184514 246174 185134 305618
rect 184514 245938 184546 246174
rect 184782 245938 184866 246174
rect 185102 245938 185134 246174
rect 184514 245854 185134 245938
rect 184514 245618 184546 245854
rect 184782 245618 184866 245854
rect 185102 245618 185134 245854
rect 184514 186174 185134 245618
rect 184514 185938 184546 186174
rect 184782 185938 184866 186174
rect 185102 185938 185134 186174
rect 184514 185854 185134 185938
rect 184514 185618 184546 185854
rect 184782 185618 184866 185854
rect 185102 185618 185134 185854
rect 184514 126174 185134 185618
rect 184514 125938 184546 126174
rect 184782 125938 184866 126174
rect 185102 125938 185134 126174
rect 184514 125854 185134 125938
rect 184514 125618 184546 125854
rect 184782 125618 184866 125854
rect 185102 125618 185134 125854
rect 184514 66174 185134 125618
rect 184514 65938 184546 66174
rect 184782 65938 184866 66174
rect 185102 65938 185134 66174
rect 184514 65854 185134 65938
rect 184514 65618 184546 65854
rect 184782 65618 184866 65854
rect 185102 65618 185134 65854
rect 184514 6174 185134 65618
rect 184514 5938 184546 6174
rect 184782 5938 184866 6174
rect 185102 5938 185134 6174
rect 184514 5854 185134 5938
rect 184514 5618 184546 5854
rect 184782 5618 184866 5854
rect 185102 5618 185134 5854
rect 184514 -2266 185134 5618
rect 184514 -2502 184546 -2266
rect 184782 -2502 184866 -2266
rect 185102 -2502 185134 -2266
rect 184514 -2586 185134 -2502
rect 184514 -2822 184546 -2586
rect 184782 -2822 184866 -2586
rect 185102 -2822 185134 -2586
rect 184514 -3814 185134 -2822
rect 188234 669894 188854 708122
rect 188234 669658 188266 669894
rect 188502 669658 188586 669894
rect 188822 669658 188854 669894
rect 188234 669574 188854 669658
rect 188234 669338 188266 669574
rect 188502 669338 188586 669574
rect 188822 669338 188854 669574
rect 188234 609894 188854 669338
rect 188234 609658 188266 609894
rect 188502 609658 188586 609894
rect 188822 609658 188854 609894
rect 188234 609574 188854 609658
rect 188234 609338 188266 609574
rect 188502 609338 188586 609574
rect 188822 609338 188854 609574
rect 188234 549894 188854 609338
rect 188234 549658 188266 549894
rect 188502 549658 188586 549894
rect 188822 549658 188854 549894
rect 188234 549574 188854 549658
rect 188234 549338 188266 549574
rect 188502 549338 188586 549574
rect 188822 549338 188854 549574
rect 188234 489894 188854 549338
rect 188234 489658 188266 489894
rect 188502 489658 188586 489894
rect 188822 489658 188854 489894
rect 188234 489574 188854 489658
rect 188234 489338 188266 489574
rect 188502 489338 188586 489574
rect 188822 489338 188854 489574
rect 188234 429894 188854 489338
rect 188234 429658 188266 429894
rect 188502 429658 188586 429894
rect 188822 429658 188854 429894
rect 188234 429574 188854 429658
rect 188234 429338 188266 429574
rect 188502 429338 188586 429574
rect 188822 429338 188854 429574
rect 188234 369894 188854 429338
rect 188234 369658 188266 369894
rect 188502 369658 188586 369894
rect 188822 369658 188854 369894
rect 188234 369574 188854 369658
rect 188234 369338 188266 369574
rect 188502 369338 188586 369574
rect 188822 369338 188854 369574
rect 188234 309894 188854 369338
rect 188234 309658 188266 309894
rect 188502 309658 188586 309894
rect 188822 309658 188854 309894
rect 188234 309574 188854 309658
rect 188234 309338 188266 309574
rect 188502 309338 188586 309574
rect 188822 309338 188854 309574
rect 188234 249894 188854 309338
rect 188234 249658 188266 249894
rect 188502 249658 188586 249894
rect 188822 249658 188854 249894
rect 188234 249574 188854 249658
rect 188234 249338 188266 249574
rect 188502 249338 188586 249574
rect 188822 249338 188854 249574
rect 188234 189894 188854 249338
rect 188234 189658 188266 189894
rect 188502 189658 188586 189894
rect 188822 189658 188854 189894
rect 188234 189574 188854 189658
rect 188234 189338 188266 189574
rect 188502 189338 188586 189574
rect 188822 189338 188854 189574
rect 188234 129894 188854 189338
rect 188234 129658 188266 129894
rect 188502 129658 188586 129894
rect 188822 129658 188854 129894
rect 188234 129574 188854 129658
rect 188234 129338 188266 129574
rect 188502 129338 188586 129574
rect 188822 129338 188854 129574
rect 188234 69894 188854 129338
rect 188234 69658 188266 69894
rect 188502 69658 188586 69894
rect 188822 69658 188854 69894
rect 188234 69574 188854 69658
rect 188234 69338 188266 69574
rect 188502 69338 188586 69574
rect 188822 69338 188854 69574
rect 188234 9894 188854 69338
rect 188234 9658 188266 9894
rect 188502 9658 188586 9894
rect 188822 9658 188854 9894
rect 188234 9574 188854 9658
rect 188234 9338 188266 9574
rect 188502 9338 188586 9574
rect 188822 9338 188854 9574
rect 188234 -4186 188854 9338
rect 188234 -4422 188266 -4186
rect 188502 -4422 188586 -4186
rect 188822 -4422 188854 -4186
rect 188234 -4506 188854 -4422
rect 188234 -4742 188266 -4506
rect 188502 -4742 188586 -4506
rect 188822 -4742 188854 -4506
rect 188234 -5734 188854 -4742
rect 191954 673614 192574 710042
rect 221954 711558 222574 711590
rect 221954 711322 221986 711558
rect 222222 711322 222306 711558
rect 222542 711322 222574 711558
rect 221954 711238 222574 711322
rect 221954 711002 221986 711238
rect 222222 711002 222306 711238
rect 222542 711002 222574 711238
rect 218234 709638 218854 709670
rect 218234 709402 218266 709638
rect 218502 709402 218586 709638
rect 218822 709402 218854 709638
rect 218234 709318 218854 709402
rect 218234 709082 218266 709318
rect 218502 709082 218586 709318
rect 218822 709082 218854 709318
rect 214514 707718 215134 707750
rect 214514 707482 214546 707718
rect 214782 707482 214866 707718
rect 215102 707482 215134 707718
rect 214514 707398 215134 707482
rect 214514 707162 214546 707398
rect 214782 707162 214866 707398
rect 215102 707162 215134 707398
rect 191954 673378 191986 673614
rect 192222 673378 192306 673614
rect 192542 673378 192574 673614
rect 191954 673294 192574 673378
rect 191954 673058 191986 673294
rect 192222 673058 192306 673294
rect 192542 673058 192574 673294
rect 191954 613614 192574 673058
rect 191954 613378 191986 613614
rect 192222 613378 192306 613614
rect 192542 613378 192574 613614
rect 191954 613294 192574 613378
rect 191954 613058 191986 613294
rect 192222 613058 192306 613294
rect 192542 613058 192574 613294
rect 191954 553614 192574 613058
rect 191954 553378 191986 553614
rect 192222 553378 192306 553614
rect 192542 553378 192574 553614
rect 191954 553294 192574 553378
rect 191954 553058 191986 553294
rect 192222 553058 192306 553294
rect 192542 553058 192574 553294
rect 191954 493614 192574 553058
rect 191954 493378 191986 493614
rect 192222 493378 192306 493614
rect 192542 493378 192574 493614
rect 191954 493294 192574 493378
rect 191954 493058 191986 493294
rect 192222 493058 192306 493294
rect 192542 493058 192574 493294
rect 191954 433614 192574 493058
rect 191954 433378 191986 433614
rect 192222 433378 192306 433614
rect 192542 433378 192574 433614
rect 191954 433294 192574 433378
rect 191954 433058 191986 433294
rect 192222 433058 192306 433294
rect 192542 433058 192574 433294
rect 191954 373614 192574 433058
rect 191954 373378 191986 373614
rect 192222 373378 192306 373614
rect 192542 373378 192574 373614
rect 191954 373294 192574 373378
rect 191954 373058 191986 373294
rect 192222 373058 192306 373294
rect 192542 373058 192574 373294
rect 191954 313614 192574 373058
rect 191954 313378 191986 313614
rect 192222 313378 192306 313614
rect 192542 313378 192574 313614
rect 191954 313294 192574 313378
rect 191954 313058 191986 313294
rect 192222 313058 192306 313294
rect 192542 313058 192574 313294
rect 191954 253614 192574 313058
rect 210794 705798 211414 705830
rect 210794 705562 210826 705798
rect 211062 705562 211146 705798
rect 211382 705562 211414 705798
rect 210794 705478 211414 705562
rect 210794 705242 210826 705478
rect 211062 705242 211146 705478
rect 211382 705242 211414 705478
rect 210794 692454 211414 705242
rect 210794 692218 210826 692454
rect 211062 692218 211146 692454
rect 211382 692218 211414 692454
rect 210794 692134 211414 692218
rect 210794 691898 210826 692134
rect 211062 691898 211146 692134
rect 211382 691898 211414 692134
rect 210794 632454 211414 691898
rect 210794 632218 210826 632454
rect 211062 632218 211146 632454
rect 211382 632218 211414 632454
rect 210794 632134 211414 632218
rect 210794 631898 210826 632134
rect 211062 631898 211146 632134
rect 211382 631898 211414 632134
rect 210794 572454 211414 631898
rect 210794 572218 210826 572454
rect 211062 572218 211146 572454
rect 211382 572218 211414 572454
rect 210794 572134 211414 572218
rect 210794 571898 210826 572134
rect 211062 571898 211146 572134
rect 211382 571898 211414 572134
rect 210794 512454 211414 571898
rect 210794 512218 210826 512454
rect 211062 512218 211146 512454
rect 211382 512218 211414 512454
rect 210794 512134 211414 512218
rect 210794 511898 210826 512134
rect 211062 511898 211146 512134
rect 211382 511898 211414 512134
rect 210794 452454 211414 511898
rect 210794 452218 210826 452454
rect 211062 452218 211146 452454
rect 211382 452218 211414 452454
rect 210794 452134 211414 452218
rect 210794 451898 210826 452134
rect 211062 451898 211146 452134
rect 211382 451898 211414 452134
rect 210794 392454 211414 451898
rect 210794 392218 210826 392454
rect 211062 392218 211146 392454
rect 211382 392218 211414 392454
rect 210794 392134 211414 392218
rect 210794 391898 210826 392134
rect 211062 391898 211146 392134
rect 211382 391898 211414 392134
rect 210794 332454 211414 391898
rect 210794 332218 210826 332454
rect 211062 332218 211146 332454
rect 211382 332218 211414 332454
rect 210794 332134 211414 332218
rect 210794 331898 210826 332134
rect 211062 331898 211146 332134
rect 211382 331898 211414 332134
rect 210794 272454 211414 331898
rect 210794 272218 210826 272454
rect 211062 272218 211146 272454
rect 211382 272218 211414 272454
rect 210794 272134 211414 272218
rect 210794 271898 210826 272134
rect 211062 271898 211146 272134
rect 211382 271898 211414 272134
rect 210794 254295 211414 271898
rect 214514 696174 215134 707162
rect 214514 695938 214546 696174
rect 214782 695938 214866 696174
rect 215102 695938 215134 696174
rect 214514 695854 215134 695938
rect 214514 695618 214546 695854
rect 214782 695618 214866 695854
rect 215102 695618 215134 695854
rect 214514 636174 215134 695618
rect 214514 635938 214546 636174
rect 214782 635938 214866 636174
rect 215102 635938 215134 636174
rect 214514 635854 215134 635938
rect 214514 635618 214546 635854
rect 214782 635618 214866 635854
rect 215102 635618 215134 635854
rect 214514 576174 215134 635618
rect 214514 575938 214546 576174
rect 214782 575938 214866 576174
rect 215102 575938 215134 576174
rect 214514 575854 215134 575938
rect 214514 575618 214546 575854
rect 214782 575618 214866 575854
rect 215102 575618 215134 575854
rect 214514 516174 215134 575618
rect 214514 515938 214546 516174
rect 214782 515938 214866 516174
rect 215102 515938 215134 516174
rect 214514 515854 215134 515938
rect 214514 515618 214546 515854
rect 214782 515618 214866 515854
rect 215102 515618 215134 515854
rect 214514 456174 215134 515618
rect 214514 455938 214546 456174
rect 214782 455938 214866 456174
rect 215102 455938 215134 456174
rect 214514 455854 215134 455938
rect 214514 455618 214546 455854
rect 214782 455618 214866 455854
rect 215102 455618 215134 455854
rect 214514 396174 215134 455618
rect 214514 395938 214546 396174
rect 214782 395938 214866 396174
rect 215102 395938 215134 396174
rect 214514 395854 215134 395938
rect 214514 395618 214546 395854
rect 214782 395618 214866 395854
rect 215102 395618 215134 395854
rect 214514 336174 215134 395618
rect 214514 335938 214546 336174
rect 214782 335938 214866 336174
rect 215102 335938 215134 336174
rect 214514 335854 215134 335938
rect 214514 335618 214546 335854
rect 214782 335618 214866 335854
rect 215102 335618 215134 335854
rect 214514 276174 215134 335618
rect 214514 275938 214546 276174
rect 214782 275938 214866 276174
rect 215102 275938 215134 276174
rect 214514 275854 215134 275938
rect 214514 275618 214546 275854
rect 214782 275618 214866 275854
rect 215102 275618 215134 275854
rect 214514 254295 215134 275618
rect 218234 699894 218854 709082
rect 218234 699658 218266 699894
rect 218502 699658 218586 699894
rect 218822 699658 218854 699894
rect 219203 699820 219269 699821
rect 219203 699756 219204 699820
rect 219268 699756 219269 699820
rect 219203 699755 219269 699756
rect 218234 699574 218854 699658
rect 218234 699338 218266 699574
rect 218502 699338 218586 699574
rect 218822 699338 218854 699574
rect 218234 639894 218854 699338
rect 218234 639658 218266 639894
rect 218502 639658 218586 639894
rect 218822 639658 218854 639894
rect 218234 639574 218854 639658
rect 218234 639338 218266 639574
rect 218502 639338 218586 639574
rect 218822 639338 218854 639574
rect 218234 579894 218854 639338
rect 218234 579658 218266 579894
rect 218502 579658 218586 579894
rect 218822 579658 218854 579894
rect 218234 579574 218854 579658
rect 218234 579338 218266 579574
rect 218502 579338 218586 579574
rect 218822 579338 218854 579574
rect 218234 519894 218854 579338
rect 218234 519658 218266 519894
rect 218502 519658 218586 519894
rect 218822 519658 218854 519894
rect 218234 519574 218854 519658
rect 218234 519338 218266 519574
rect 218502 519338 218586 519574
rect 218822 519338 218854 519574
rect 218234 459894 218854 519338
rect 218234 459658 218266 459894
rect 218502 459658 218586 459894
rect 218822 459658 218854 459894
rect 218234 459574 218854 459658
rect 218234 459338 218266 459574
rect 218502 459338 218586 459574
rect 218822 459338 218854 459574
rect 218234 399894 218854 459338
rect 218234 399658 218266 399894
rect 218502 399658 218586 399894
rect 218822 399658 218854 399894
rect 218234 399574 218854 399658
rect 218234 399338 218266 399574
rect 218502 399338 218586 399574
rect 218822 399338 218854 399574
rect 218234 339894 218854 399338
rect 218234 339658 218266 339894
rect 218502 339658 218586 339894
rect 218822 339658 218854 339894
rect 218234 339574 218854 339658
rect 218234 339338 218266 339574
rect 218502 339338 218586 339574
rect 218822 339338 218854 339574
rect 218234 279894 218854 339338
rect 218234 279658 218266 279894
rect 218502 279658 218586 279894
rect 218822 279658 218854 279894
rect 218234 279574 218854 279658
rect 218234 279338 218266 279574
rect 218502 279338 218586 279574
rect 218822 279338 218854 279574
rect 218234 254295 218854 279338
rect 191954 253378 191986 253614
rect 192222 253378 192306 253614
rect 192542 253378 192574 253614
rect 191954 253294 192574 253378
rect 191954 253058 191986 253294
rect 192222 253058 192306 253294
rect 192542 253058 192574 253294
rect 191954 193614 192574 253058
rect 210555 251700 210621 251701
rect 210555 251636 210556 251700
rect 210620 251636 210621 251700
rect 210555 251635 210621 251636
rect 204208 242454 204528 242486
rect 204208 242218 204250 242454
rect 204486 242218 204528 242454
rect 204208 242134 204528 242218
rect 204208 241898 204250 242134
rect 204486 241898 204528 242134
rect 204208 241866 204528 241898
rect 191954 193378 191986 193614
rect 192222 193378 192306 193614
rect 192542 193378 192574 193614
rect 191954 193294 192574 193378
rect 191954 193058 191986 193294
rect 192222 193058 192306 193294
rect 192542 193058 192574 193294
rect 191954 133614 192574 193058
rect 191954 133378 191986 133614
rect 192222 133378 192306 133614
rect 192542 133378 192574 133614
rect 191954 133294 192574 133378
rect 191954 133058 191986 133294
rect 192222 133058 192306 133294
rect 192542 133058 192574 133294
rect 191954 73614 192574 133058
rect 191954 73378 191986 73614
rect 192222 73378 192306 73614
rect 192542 73378 192574 73614
rect 191954 73294 192574 73378
rect 191954 73058 191986 73294
rect 192222 73058 192306 73294
rect 192542 73058 192574 73294
rect 191954 13614 192574 73058
rect 191954 13378 191986 13614
rect 192222 13378 192306 13614
rect 192542 13378 192574 13614
rect 191954 13294 192574 13378
rect 191954 13058 191986 13294
rect 192222 13058 192306 13294
rect 192542 13058 192574 13294
rect 161954 -7302 161986 -7066
rect 162222 -7302 162306 -7066
rect 162542 -7302 162574 -7066
rect 161954 -7386 162574 -7302
rect 161954 -7622 161986 -7386
rect 162222 -7622 162306 -7386
rect 162542 -7622 162574 -7386
rect 161954 -7654 162574 -7622
rect 191954 -6106 192574 13058
rect 210558 5677 210618 251635
rect 219206 238770 219266 699755
rect 221954 643614 222574 711002
rect 251954 710598 252574 711590
rect 251954 710362 251986 710598
rect 252222 710362 252306 710598
rect 252542 710362 252574 710598
rect 251954 710278 252574 710362
rect 251954 710042 251986 710278
rect 252222 710042 252306 710278
rect 252542 710042 252574 710278
rect 248234 708678 248854 709670
rect 248234 708442 248266 708678
rect 248502 708442 248586 708678
rect 248822 708442 248854 708678
rect 248234 708358 248854 708442
rect 248234 708122 248266 708358
rect 248502 708122 248586 708358
rect 248822 708122 248854 708358
rect 244514 706758 245134 707750
rect 244514 706522 244546 706758
rect 244782 706522 244866 706758
rect 245102 706522 245134 706758
rect 244514 706438 245134 706522
rect 244514 706202 244546 706438
rect 244782 706202 244866 706438
rect 245102 706202 245134 706438
rect 221954 643378 221986 643614
rect 222222 643378 222306 643614
rect 222542 643378 222574 643614
rect 221954 643294 222574 643378
rect 221954 643058 221986 643294
rect 222222 643058 222306 643294
rect 222542 643058 222574 643294
rect 221954 583614 222574 643058
rect 221954 583378 221986 583614
rect 222222 583378 222306 583614
rect 222542 583378 222574 583614
rect 221954 583294 222574 583378
rect 221954 583058 221986 583294
rect 222222 583058 222306 583294
rect 222542 583058 222574 583294
rect 221954 523614 222574 583058
rect 221954 523378 221986 523614
rect 222222 523378 222306 523614
rect 222542 523378 222574 523614
rect 221954 523294 222574 523378
rect 221954 523058 221986 523294
rect 222222 523058 222306 523294
rect 222542 523058 222574 523294
rect 221954 463614 222574 523058
rect 221954 463378 221986 463614
rect 222222 463378 222306 463614
rect 222542 463378 222574 463614
rect 221954 463294 222574 463378
rect 221954 463058 221986 463294
rect 222222 463058 222306 463294
rect 222542 463058 222574 463294
rect 221954 403614 222574 463058
rect 221954 403378 221986 403614
rect 222222 403378 222306 403614
rect 222542 403378 222574 403614
rect 221954 403294 222574 403378
rect 221954 403058 221986 403294
rect 222222 403058 222306 403294
rect 222542 403058 222574 403294
rect 221954 343614 222574 403058
rect 221954 343378 221986 343614
rect 222222 343378 222306 343614
rect 222542 343378 222574 343614
rect 221954 343294 222574 343378
rect 221954 343058 221986 343294
rect 222222 343058 222306 343294
rect 222542 343058 222574 343294
rect 221954 283614 222574 343058
rect 221954 283378 221986 283614
rect 222222 283378 222306 283614
rect 222542 283378 222574 283614
rect 221954 283294 222574 283378
rect 221954 283058 221986 283294
rect 222222 283058 222306 283294
rect 222542 283058 222574 283294
rect 221954 254295 222574 283058
rect 240794 704838 241414 705830
rect 240794 704602 240826 704838
rect 241062 704602 241146 704838
rect 241382 704602 241414 704838
rect 240794 704518 241414 704602
rect 240794 704282 240826 704518
rect 241062 704282 241146 704518
rect 241382 704282 241414 704518
rect 240794 662454 241414 704282
rect 240794 662218 240826 662454
rect 241062 662218 241146 662454
rect 241382 662218 241414 662454
rect 240794 662134 241414 662218
rect 240794 661898 240826 662134
rect 241062 661898 241146 662134
rect 241382 661898 241414 662134
rect 240794 602454 241414 661898
rect 240794 602218 240826 602454
rect 241062 602218 241146 602454
rect 241382 602218 241414 602454
rect 240794 602134 241414 602218
rect 240794 601898 240826 602134
rect 241062 601898 241146 602134
rect 241382 601898 241414 602134
rect 240794 542454 241414 601898
rect 240794 542218 240826 542454
rect 241062 542218 241146 542454
rect 241382 542218 241414 542454
rect 240794 542134 241414 542218
rect 240794 541898 240826 542134
rect 241062 541898 241146 542134
rect 241382 541898 241414 542134
rect 240794 482454 241414 541898
rect 240794 482218 240826 482454
rect 241062 482218 241146 482454
rect 241382 482218 241414 482454
rect 240794 482134 241414 482218
rect 240794 481898 240826 482134
rect 241062 481898 241146 482134
rect 241382 481898 241414 482134
rect 240794 422454 241414 481898
rect 240794 422218 240826 422454
rect 241062 422218 241146 422454
rect 241382 422218 241414 422454
rect 240794 422134 241414 422218
rect 240794 421898 240826 422134
rect 241062 421898 241146 422134
rect 241382 421898 241414 422134
rect 240794 362454 241414 421898
rect 240794 362218 240826 362454
rect 241062 362218 241146 362454
rect 241382 362218 241414 362454
rect 240794 362134 241414 362218
rect 240794 361898 240826 362134
rect 241062 361898 241146 362134
rect 241382 361898 241414 362134
rect 240794 302454 241414 361898
rect 240794 302218 240826 302454
rect 241062 302218 241146 302454
rect 241382 302218 241414 302454
rect 240794 302134 241414 302218
rect 240794 301898 240826 302134
rect 241062 301898 241146 302134
rect 241382 301898 241414 302134
rect 240794 254295 241414 301898
rect 244514 666174 245134 706202
rect 244514 665938 244546 666174
rect 244782 665938 244866 666174
rect 245102 665938 245134 666174
rect 244514 665854 245134 665938
rect 244514 665618 244546 665854
rect 244782 665618 244866 665854
rect 245102 665618 245134 665854
rect 244514 606174 245134 665618
rect 244514 605938 244546 606174
rect 244782 605938 244866 606174
rect 245102 605938 245134 606174
rect 244514 605854 245134 605938
rect 244514 605618 244546 605854
rect 244782 605618 244866 605854
rect 245102 605618 245134 605854
rect 244514 546174 245134 605618
rect 244514 545938 244546 546174
rect 244782 545938 244866 546174
rect 245102 545938 245134 546174
rect 244514 545854 245134 545938
rect 244514 545618 244546 545854
rect 244782 545618 244866 545854
rect 245102 545618 245134 545854
rect 244514 486174 245134 545618
rect 244514 485938 244546 486174
rect 244782 485938 244866 486174
rect 245102 485938 245134 486174
rect 244514 485854 245134 485938
rect 244514 485618 244546 485854
rect 244782 485618 244866 485854
rect 245102 485618 245134 485854
rect 244514 426174 245134 485618
rect 244514 425938 244546 426174
rect 244782 425938 244866 426174
rect 245102 425938 245134 426174
rect 244514 425854 245134 425938
rect 244514 425618 244546 425854
rect 244782 425618 244866 425854
rect 245102 425618 245134 425854
rect 244514 366174 245134 425618
rect 244514 365938 244546 366174
rect 244782 365938 244866 366174
rect 245102 365938 245134 366174
rect 244514 365854 245134 365938
rect 244514 365618 244546 365854
rect 244782 365618 244866 365854
rect 245102 365618 245134 365854
rect 244514 306174 245134 365618
rect 244514 305938 244546 306174
rect 244782 305938 244866 306174
rect 245102 305938 245134 306174
rect 244514 305854 245134 305938
rect 244514 305618 244546 305854
rect 244782 305618 244866 305854
rect 245102 305618 245134 305854
rect 244514 254295 245134 305618
rect 248234 669894 248854 708122
rect 248234 669658 248266 669894
rect 248502 669658 248586 669894
rect 248822 669658 248854 669894
rect 248234 669574 248854 669658
rect 248234 669338 248266 669574
rect 248502 669338 248586 669574
rect 248822 669338 248854 669574
rect 248234 609894 248854 669338
rect 248234 609658 248266 609894
rect 248502 609658 248586 609894
rect 248822 609658 248854 609894
rect 248234 609574 248854 609658
rect 248234 609338 248266 609574
rect 248502 609338 248586 609574
rect 248822 609338 248854 609574
rect 248234 549894 248854 609338
rect 248234 549658 248266 549894
rect 248502 549658 248586 549894
rect 248822 549658 248854 549894
rect 248234 549574 248854 549658
rect 248234 549338 248266 549574
rect 248502 549338 248586 549574
rect 248822 549338 248854 549574
rect 248234 489894 248854 549338
rect 248234 489658 248266 489894
rect 248502 489658 248586 489894
rect 248822 489658 248854 489894
rect 248234 489574 248854 489658
rect 248234 489338 248266 489574
rect 248502 489338 248586 489574
rect 248822 489338 248854 489574
rect 248234 429894 248854 489338
rect 248234 429658 248266 429894
rect 248502 429658 248586 429894
rect 248822 429658 248854 429894
rect 248234 429574 248854 429658
rect 248234 429338 248266 429574
rect 248502 429338 248586 429574
rect 248822 429338 248854 429574
rect 248234 369894 248854 429338
rect 248234 369658 248266 369894
rect 248502 369658 248586 369894
rect 248822 369658 248854 369894
rect 248234 369574 248854 369658
rect 248234 369338 248266 369574
rect 248502 369338 248586 369574
rect 248822 369338 248854 369574
rect 248234 309894 248854 369338
rect 248234 309658 248266 309894
rect 248502 309658 248586 309894
rect 248822 309658 248854 309894
rect 248234 309574 248854 309658
rect 248234 309338 248266 309574
rect 248502 309338 248586 309574
rect 248822 309338 248854 309574
rect 248234 254295 248854 309338
rect 251954 673614 252574 710042
rect 281954 711558 282574 711590
rect 281954 711322 281986 711558
rect 282222 711322 282306 711558
rect 282542 711322 282574 711558
rect 281954 711238 282574 711322
rect 281954 711002 281986 711238
rect 282222 711002 282306 711238
rect 282542 711002 282574 711238
rect 278234 709638 278854 709670
rect 278234 709402 278266 709638
rect 278502 709402 278586 709638
rect 278822 709402 278854 709638
rect 278234 709318 278854 709402
rect 278234 709082 278266 709318
rect 278502 709082 278586 709318
rect 278822 709082 278854 709318
rect 274514 707718 275134 707750
rect 274514 707482 274546 707718
rect 274782 707482 274866 707718
rect 275102 707482 275134 707718
rect 274514 707398 275134 707482
rect 274514 707162 274546 707398
rect 274782 707162 274866 707398
rect 275102 707162 275134 707398
rect 251954 673378 251986 673614
rect 252222 673378 252306 673614
rect 252542 673378 252574 673614
rect 251954 673294 252574 673378
rect 251954 673058 251986 673294
rect 252222 673058 252306 673294
rect 252542 673058 252574 673294
rect 251954 613614 252574 673058
rect 251954 613378 251986 613614
rect 252222 613378 252306 613614
rect 252542 613378 252574 613614
rect 251954 613294 252574 613378
rect 251954 613058 251986 613294
rect 252222 613058 252306 613294
rect 252542 613058 252574 613294
rect 251954 553614 252574 613058
rect 251954 553378 251986 553614
rect 252222 553378 252306 553614
rect 252542 553378 252574 553614
rect 251954 553294 252574 553378
rect 251954 553058 251986 553294
rect 252222 553058 252306 553294
rect 252542 553058 252574 553294
rect 251954 493614 252574 553058
rect 251954 493378 251986 493614
rect 252222 493378 252306 493614
rect 252542 493378 252574 493614
rect 251954 493294 252574 493378
rect 251954 493058 251986 493294
rect 252222 493058 252306 493294
rect 252542 493058 252574 493294
rect 251954 433614 252574 493058
rect 251954 433378 251986 433614
rect 252222 433378 252306 433614
rect 252542 433378 252574 433614
rect 251954 433294 252574 433378
rect 251954 433058 251986 433294
rect 252222 433058 252306 433294
rect 252542 433058 252574 433294
rect 251954 373614 252574 433058
rect 251954 373378 251986 373614
rect 252222 373378 252306 373614
rect 252542 373378 252574 373614
rect 251954 373294 252574 373378
rect 251954 373058 251986 373294
rect 252222 373058 252306 373294
rect 252542 373058 252574 373294
rect 251954 313614 252574 373058
rect 251954 313378 251986 313614
rect 252222 313378 252306 313614
rect 252542 313378 252574 313614
rect 251954 313294 252574 313378
rect 251954 313058 251986 313294
rect 252222 313058 252306 313294
rect 252542 313058 252574 313294
rect 251954 254295 252574 313058
rect 270794 705798 271414 705830
rect 270794 705562 270826 705798
rect 271062 705562 271146 705798
rect 271382 705562 271414 705798
rect 270794 705478 271414 705562
rect 270794 705242 270826 705478
rect 271062 705242 271146 705478
rect 271382 705242 271414 705478
rect 270794 692454 271414 705242
rect 270794 692218 270826 692454
rect 271062 692218 271146 692454
rect 271382 692218 271414 692454
rect 270794 692134 271414 692218
rect 270794 691898 270826 692134
rect 271062 691898 271146 692134
rect 271382 691898 271414 692134
rect 270794 632454 271414 691898
rect 270794 632218 270826 632454
rect 271062 632218 271146 632454
rect 271382 632218 271414 632454
rect 270794 632134 271414 632218
rect 270794 631898 270826 632134
rect 271062 631898 271146 632134
rect 271382 631898 271414 632134
rect 270794 572454 271414 631898
rect 270794 572218 270826 572454
rect 271062 572218 271146 572454
rect 271382 572218 271414 572454
rect 270794 572134 271414 572218
rect 270794 571898 270826 572134
rect 271062 571898 271146 572134
rect 271382 571898 271414 572134
rect 270794 512454 271414 571898
rect 270794 512218 270826 512454
rect 271062 512218 271146 512454
rect 271382 512218 271414 512454
rect 270794 512134 271414 512218
rect 270794 511898 270826 512134
rect 271062 511898 271146 512134
rect 271382 511898 271414 512134
rect 270794 452454 271414 511898
rect 270794 452218 270826 452454
rect 271062 452218 271146 452454
rect 271382 452218 271414 452454
rect 270794 452134 271414 452218
rect 270794 451898 270826 452134
rect 271062 451898 271146 452134
rect 271382 451898 271414 452134
rect 270794 392454 271414 451898
rect 270794 392218 270826 392454
rect 271062 392218 271146 392454
rect 271382 392218 271414 392454
rect 270794 392134 271414 392218
rect 270794 391898 270826 392134
rect 271062 391898 271146 392134
rect 271382 391898 271414 392134
rect 270794 332454 271414 391898
rect 270794 332218 270826 332454
rect 271062 332218 271146 332454
rect 271382 332218 271414 332454
rect 270794 332134 271414 332218
rect 270794 331898 270826 332134
rect 271062 331898 271146 332134
rect 271382 331898 271414 332134
rect 270794 272454 271414 331898
rect 270794 272218 270826 272454
rect 271062 272218 271146 272454
rect 271382 272218 271414 272454
rect 270794 272134 271414 272218
rect 270794 271898 270826 272134
rect 271062 271898 271146 272134
rect 271382 271898 271414 272134
rect 249566 246941 249626 247062
rect 249563 246940 249629 246941
rect 249563 246876 249564 246940
rect 249628 246876 249629 246940
rect 249563 246875 249629 246876
rect 234928 242454 235248 242486
rect 234928 242218 234970 242454
rect 235206 242218 235248 242454
rect 234928 242134 235248 242218
rect 234928 241898 234970 242134
rect 235206 241898 235248 242134
rect 234928 241866 235248 241898
rect 218286 238710 219266 238770
rect 218286 218058 218346 238710
rect 249566 217701 249626 217822
rect 249563 217700 249629 217701
rect 249563 217636 249564 217700
rect 249628 217636 249629 217700
rect 249563 217635 249629 217636
rect 219568 212454 219888 212486
rect 219568 212218 219610 212454
rect 219846 212218 219888 212454
rect 219568 212134 219888 212218
rect 219568 211898 219610 212134
rect 219846 211898 219888 212134
rect 219568 211866 219888 211898
rect 270794 212454 271414 271898
rect 270794 212218 270826 212454
rect 271062 212218 271146 212454
rect 271382 212218 271414 212454
rect 270794 212134 271414 212218
rect 270794 211898 270826 212134
rect 271062 211898 271146 212134
rect 271382 211898 271414 212134
rect 249563 205052 249629 205053
rect 249563 204988 249564 205052
rect 249628 204988 249629 205052
rect 249563 204987 249629 204988
rect 249566 204458 249626 204987
rect 210794 152454 211414 198000
rect 210794 152218 210826 152454
rect 211062 152218 211146 152454
rect 211382 152218 211414 152454
rect 210794 152134 211414 152218
rect 210794 151898 210826 152134
rect 211062 151898 211146 152134
rect 211382 151898 211414 152134
rect 210794 92454 211414 151898
rect 210794 92218 210826 92454
rect 211062 92218 211146 92454
rect 211382 92218 211414 92454
rect 210794 92134 211414 92218
rect 210794 91898 210826 92134
rect 211062 91898 211146 92134
rect 211382 91898 211414 92134
rect 210794 32454 211414 91898
rect 210794 32218 210826 32454
rect 211062 32218 211146 32454
rect 211382 32218 211414 32454
rect 210794 32134 211414 32218
rect 210794 31898 210826 32134
rect 211062 31898 211146 32134
rect 211382 31898 211414 32134
rect 210555 5676 210621 5677
rect 210555 5612 210556 5676
rect 210620 5612 210621 5676
rect 210555 5611 210621 5612
rect 210794 -1306 211414 31898
rect 210794 -1542 210826 -1306
rect 211062 -1542 211146 -1306
rect 211382 -1542 211414 -1306
rect 210794 -1626 211414 -1542
rect 210794 -1862 210826 -1626
rect 211062 -1862 211146 -1626
rect 211382 -1862 211414 -1626
rect 210794 -1894 211414 -1862
rect 214514 156174 215134 198000
rect 214514 155938 214546 156174
rect 214782 155938 214866 156174
rect 215102 155938 215134 156174
rect 214514 155854 215134 155938
rect 214514 155618 214546 155854
rect 214782 155618 214866 155854
rect 215102 155618 215134 155854
rect 214514 96174 215134 155618
rect 214514 95938 214546 96174
rect 214782 95938 214866 96174
rect 215102 95938 215134 96174
rect 214514 95854 215134 95938
rect 214514 95618 214546 95854
rect 214782 95618 214866 95854
rect 215102 95618 215134 95854
rect 214514 36174 215134 95618
rect 214514 35938 214546 36174
rect 214782 35938 214866 36174
rect 215102 35938 215134 36174
rect 214514 35854 215134 35938
rect 214514 35618 214546 35854
rect 214782 35618 214866 35854
rect 215102 35618 215134 35854
rect 214514 -3226 215134 35618
rect 214514 -3462 214546 -3226
rect 214782 -3462 214866 -3226
rect 215102 -3462 215134 -3226
rect 214514 -3546 215134 -3462
rect 214514 -3782 214546 -3546
rect 214782 -3782 214866 -3546
rect 215102 -3782 215134 -3546
rect 214514 -3814 215134 -3782
rect 218234 159894 218854 198000
rect 218234 159658 218266 159894
rect 218502 159658 218586 159894
rect 218822 159658 218854 159894
rect 218234 159574 218854 159658
rect 218234 159338 218266 159574
rect 218502 159338 218586 159574
rect 218822 159338 218854 159574
rect 218234 99894 218854 159338
rect 218234 99658 218266 99894
rect 218502 99658 218586 99894
rect 218822 99658 218854 99894
rect 218234 99574 218854 99658
rect 218234 99338 218266 99574
rect 218502 99338 218586 99574
rect 218822 99338 218854 99574
rect 218234 39894 218854 99338
rect 218234 39658 218266 39894
rect 218502 39658 218586 39894
rect 218822 39658 218854 39894
rect 218234 39574 218854 39658
rect 218234 39338 218266 39574
rect 218502 39338 218586 39574
rect 218822 39338 218854 39574
rect 218234 -5146 218854 39338
rect 218234 -5382 218266 -5146
rect 218502 -5382 218586 -5146
rect 218822 -5382 218854 -5146
rect 218234 -5466 218854 -5382
rect 218234 -5702 218266 -5466
rect 218502 -5702 218586 -5466
rect 218822 -5702 218854 -5466
rect 218234 -5734 218854 -5702
rect 221954 163614 222574 198000
rect 221954 163378 221986 163614
rect 222222 163378 222306 163614
rect 222542 163378 222574 163614
rect 221954 163294 222574 163378
rect 221954 163058 221986 163294
rect 222222 163058 222306 163294
rect 222542 163058 222574 163294
rect 221954 103614 222574 163058
rect 221954 103378 221986 103614
rect 222222 103378 222306 103614
rect 222542 103378 222574 103614
rect 221954 103294 222574 103378
rect 221954 103058 221986 103294
rect 222222 103058 222306 103294
rect 222542 103058 222574 103294
rect 221954 43614 222574 103058
rect 221954 43378 221986 43614
rect 222222 43378 222306 43614
rect 222542 43378 222574 43614
rect 221954 43294 222574 43378
rect 221954 43058 221986 43294
rect 222222 43058 222306 43294
rect 222542 43058 222574 43294
rect 191954 -6342 191986 -6106
rect 192222 -6342 192306 -6106
rect 192542 -6342 192574 -6106
rect 191954 -6426 192574 -6342
rect 191954 -6662 191986 -6426
rect 192222 -6662 192306 -6426
rect 192542 -6662 192574 -6426
rect 191954 -7654 192574 -6662
rect 221954 -7066 222574 43058
rect 240794 182454 241414 198000
rect 240794 182218 240826 182454
rect 241062 182218 241146 182454
rect 241382 182218 241414 182454
rect 240794 182134 241414 182218
rect 240794 181898 240826 182134
rect 241062 181898 241146 182134
rect 241382 181898 241414 182134
rect 240794 122454 241414 181898
rect 240794 122218 240826 122454
rect 241062 122218 241146 122454
rect 241382 122218 241414 122454
rect 240794 122134 241414 122218
rect 240794 121898 240826 122134
rect 241062 121898 241146 122134
rect 241382 121898 241414 122134
rect 240794 62454 241414 121898
rect 240794 62218 240826 62454
rect 241062 62218 241146 62454
rect 241382 62218 241414 62454
rect 240794 62134 241414 62218
rect 240794 61898 240826 62134
rect 241062 61898 241146 62134
rect 241382 61898 241414 62134
rect 240794 2454 241414 61898
rect 240794 2218 240826 2454
rect 241062 2218 241146 2454
rect 241382 2218 241414 2454
rect 240794 2134 241414 2218
rect 240794 1898 240826 2134
rect 241062 1898 241146 2134
rect 241382 1898 241414 2134
rect 240794 -346 241414 1898
rect 240794 -582 240826 -346
rect 241062 -582 241146 -346
rect 241382 -582 241414 -346
rect 240794 -666 241414 -582
rect 240794 -902 240826 -666
rect 241062 -902 241146 -666
rect 241382 -902 241414 -666
rect 240794 -1894 241414 -902
rect 244514 186174 245134 198000
rect 244514 185938 244546 186174
rect 244782 185938 244866 186174
rect 245102 185938 245134 186174
rect 244514 185854 245134 185938
rect 244514 185618 244546 185854
rect 244782 185618 244866 185854
rect 245102 185618 245134 185854
rect 244514 126174 245134 185618
rect 244514 125938 244546 126174
rect 244782 125938 244866 126174
rect 245102 125938 245134 126174
rect 244514 125854 245134 125938
rect 244514 125618 244546 125854
rect 244782 125618 244866 125854
rect 245102 125618 245134 125854
rect 244514 66174 245134 125618
rect 244514 65938 244546 66174
rect 244782 65938 244866 66174
rect 245102 65938 245134 66174
rect 244514 65854 245134 65938
rect 244514 65618 244546 65854
rect 244782 65618 244866 65854
rect 245102 65618 245134 65854
rect 244514 6174 245134 65618
rect 244514 5938 244546 6174
rect 244782 5938 244866 6174
rect 245102 5938 245134 6174
rect 244514 5854 245134 5938
rect 244514 5618 244546 5854
rect 244782 5618 244866 5854
rect 245102 5618 245134 5854
rect 244514 -2266 245134 5618
rect 244514 -2502 244546 -2266
rect 244782 -2502 244866 -2266
rect 245102 -2502 245134 -2266
rect 244514 -2586 245134 -2502
rect 244514 -2822 244546 -2586
rect 244782 -2822 244866 -2586
rect 245102 -2822 245134 -2586
rect 244514 -3814 245134 -2822
rect 248234 189894 248854 198000
rect 248234 189658 248266 189894
rect 248502 189658 248586 189894
rect 248822 189658 248854 189894
rect 248234 189574 248854 189658
rect 248234 189338 248266 189574
rect 248502 189338 248586 189574
rect 248822 189338 248854 189574
rect 248234 129894 248854 189338
rect 248234 129658 248266 129894
rect 248502 129658 248586 129894
rect 248822 129658 248854 129894
rect 248234 129574 248854 129658
rect 248234 129338 248266 129574
rect 248502 129338 248586 129574
rect 248822 129338 248854 129574
rect 248234 69894 248854 129338
rect 248234 69658 248266 69894
rect 248502 69658 248586 69894
rect 248822 69658 248854 69894
rect 248234 69574 248854 69658
rect 248234 69338 248266 69574
rect 248502 69338 248586 69574
rect 248822 69338 248854 69574
rect 248234 9894 248854 69338
rect 248234 9658 248266 9894
rect 248502 9658 248586 9894
rect 248822 9658 248854 9894
rect 248234 9574 248854 9658
rect 248234 9338 248266 9574
rect 248502 9338 248586 9574
rect 248822 9338 248854 9574
rect 248234 -4186 248854 9338
rect 248234 -4422 248266 -4186
rect 248502 -4422 248586 -4186
rect 248822 -4422 248854 -4186
rect 248234 -4506 248854 -4422
rect 248234 -4742 248266 -4506
rect 248502 -4742 248586 -4506
rect 248822 -4742 248854 -4506
rect 248234 -5734 248854 -4742
rect 251954 193614 252574 198000
rect 251954 193378 251986 193614
rect 252222 193378 252306 193614
rect 252542 193378 252574 193614
rect 251954 193294 252574 193378
rect 251954 193058 251986 193294
rect 252222 193058 252306 193294
rect 252542 193058 252574 193294
rect 251954 133614 252574 193058
rect 251954 133378 251986 133614
rect 252222 133378 252306 133614
rect 252542 133378 252574 133614
rect 251954 133294 252574 133378
rect 251954 133058 251986 133294
rect 252222 133058 252306 133294
rect 252542 133058 252574 133294
rect 251954 73614 252574 133058
rect 251954 73378 251986 73614
rect 252222 73378 252306 73614
rect 252542 73378 252574 73614
rect 251954 73294 252574 73378
rect 251954 73058 251986 73294
rect 252222 73058 252306 73294
rect 252542 73058 252574 73294
rect 251954 13614 252574 73058
rect 251954 13378 251986 13614
rect 252222 13378 252306 13614
rect 252542 13378 252574 13614
rect 251954 13294 252574 13378
rect 251954 13058 251986 13294
rect 252222 13058 252306 13294
rect 252542 13058 252574 13294
rect 221954 -7302 221986 -7066
rect 222222 -7302 222306 -7066
rect 222542 -7302 222574 -7066
rect 221954 -7386 222574 -7302
rect 221954 -7622 221986 -7386
rect 222222 -7622 222306 -7386
rect 222542 -7622 222574 -7386
rect 221954 -7654 222574 -7622
rect 251954 -6106 252574 13058
rect 270794 152454 271414 211898
rect 270794 152218 270826 152454
rect 271062 152218 271146 152454
rect 271382 152218 271414 152454
rect 270794 152134 271414 152218
rect 270794 151898 270826 152134
rect 271062 151898 271146 152134
rect 271382 151898 271414 152134
rect 270794 92454 271414 151898
rect 270794 92218 270826 92454
rect 271062 92218 271146 92454
rect 271382 92218 271414 92454
rect 270794 92134 271414 92218
rect 270794 91898 270826 92134
rect 271062 91898 271146 92134
rect 271382 91898 271414 92134
rect 270794 32454 271414 91898
rect 270794 32218 270826 32454
rect 271062 32218 271146 32454
rect 271382 32218 271414 32454
rect 270794 32134 271414 32218
rect 270794 31898 270826 32134
rect 271062 31898 271146 32134
rect 271382 31898 271414 32134
rect 270794 -1306 271414 31898
rect 270794 -1542 270826 -1306
rect 271062 -1542 271146 -1306
rect 271382 -1542 271414 -1306
rect 270794 -1626 271414 -1542
rect 270794 -1862 270826 -1626
rect 271062 -1862 271146 -1626
rect 271382 -1862 271414 -1626
rect 270794 -1894 271414 -1862
rect 274514 696174 275134 707162
rect 274514 695938 274546 696174
rect 274782 695938 274866 696174
rect 275102 695938 275134 696174
rect 274514 695854 275134 695938
rect 274514 695618 274546 695854
rect 274782 695618 274866 695854
rect 275102 695618 275134 695854
rect 274514 636174 275134 695618
rect 274514 635938 274546 636174
rect 274782 635938 274866 636174
rect 275102 635938 275134 636174
rect 274514 635854 275134 635938
rect 274514 635618 274546 635854
rect 274782 635618 274866 635854
rect 275102 635618 275134 635854
rect 274514 576174 275134 635618
rect 274514 575938 274546 576174
rect 274782 575938 274866 576174
rect 275102 575938 275134 576174
rect 274514 575854 275134 575938
rect 274514 575618 274546 575854
rect 274782 575618 274866 575854
rect 275102 575618 275134 575854
rect 274514 516174 275134 575618
rect 274514 515938 274546 516174
rect 274782 515938 274866 516174
rect 275102 515938 275134 516174
rect 274514 515854 275134 515938
rect 274514 515618 274546 515854
rect 274782 515618 274866 515854
rect 275102 515618 275134 515854
rect 274514 456174 275134 515618
rect 274514 455938 274546 456174
rect 274782 455938 274866 456174
rect 275102 455938 275134 456174
rect 274514 455854 275134 455938
rect 274514 455618 274546 455854
rect 274782 455618 274866 455854
rect 275102 455618 275134 455854
rect 274514 396174 275134 455618
rect 274514 395938 274546 396174
rect 274782 395938 274866 396174
rect 275102 395938 275134 396174
rect 274514 395854 275134 395938
rect 274514 395618 274546 395854
rect 274782 395618 274866 395854
rect 275102 395618 275134 395854
rect 274514 336174 275134 395618
rect 274514 335938 274546 336174
rect 274782 335938 274866 336174
rect 275102 335938 275134 336174
rect 274514 335854 275134 335938
rect 274514 335618 274546 335854
rect 274782 335618 274866 335854
rect 275102 335618 275134 335854
rect 274514 276174 275134 335618
rect 274514 275938 274546 276174
rect 274782 275938 274866 276174
rect 275102 275938 275134 276174
rect 274514 275854 275134 275938
rect 274514 275618 274546 275854
rect 274782 275618 274866 275854
rect 275102 275618 275134 275854
rect 274514 216174 275134 275618
rect 274514 215938 274546 216174
rect 274782 215938 274866 216174
rect 275102 215938 275134 216174
rect 274514 215854 275134 215938
rect 274514 215618 274546 215854
rect 274782 215618 274866 215854
rect 275102 215618 275134 215854
rect 274514 156174 275134 215618
rect 274514 155938 274546 156174
rect 274782 155938 274866 156174
rect 275102 155938 275134 156174
rect 274514 155854 275134 155938
rect 274514 155618 274546 155854
rect 274782 155618 274866 155854
rect 275102 155618 275134 155854
rect 274514 96174 275134 155618
rect 274514 95938 274546 96174
rect 274782 95938 274866 96174
rect 275102 95938 275134 96174
rect 274514 95854 275134 95938
rect 274514 95618 274546 95854
rect 274782 95618 274866 95854
rect 275102 95618 275134 95854
rect 274514 36174 275134 95618
rect 274514 35938 274546 36174
rect 274782 35938 274866 36174
rect 275102 35938 275134 36174
rect 274514 35854 275134 35938
rect 274514 35618 274546 35854
rect 274782 35618 274866 35854
rect 275102 35618 275134 35854
rect 274514 -3226 275134 35618
rect 274514 -3462 274546 -3226
rect 274782 -3462 274866 -3226
rect 275102 -3462 275134 -3226
rect 274514 -3546 275134 -3462
rect 274514 -3782 274546 -3546
rect 274782 -3782 274866 -3546
rect 275102 -3782 275134 -3546
rect 274514 -3814 275134 -3782
rect 278234 699894 278854 709082
rect 278234 699658 278266 699894
rect 278502 699658 278586 699894
rect 278822 699658 278854 699894
rect 278234 699574 278854 699658
rect 278234 699338 278266 699574
rect 278502 699338 278586 699574
rect 278822 699338 278854 699574
rect 278234 639894 278854 699338
rect 278234 639658 278266 639894
rect 278502 639658 278586 639894
rect 278822 639658 278854 639894
rect 278234 639574 278854 639658
rect 278234 639338 278266 639574
rect 278502 639338 278586 639574
rect 278822 639338 278854 639574
rect 278234 579894 278854 639338
rect 278234 579658 278266 579894
rect 278502 579658 278586 579894
rect 278822 579658 278854 579894
rect 278234 579574 278854 579658
rect 278234 579338 278266 579574
rect 278502 579338 278586 579574
rect 278822 579338 278854 579574
rect 278234 519894 278854 579338
rect 278234 519658 278266 519894
rect 278502 519658 278586 519894
rect 278822 519658 278854 519894
rect 278234 519574 278854 519658
rect 278234 519338 278266 519574
rect 278502 519338 278586 519574
rect 278822 519338 278854 519574
rect 278234 459894 278854 519338
rect 278234 459658 278266 459894
rect 278502 459658 278586 459894
rect 278822 459658 278854 459894
rect 278234 459574 278854 459658
rect 278234 459338 278266 459574
rect 278502 459338 278586 459574
rect 278822 459338 278854 459574
rect 278234 399894 278854 459338
rect 278234 399658 278266 399894
rect 278502 399658 278586 399894
rect 278822 399658 278854 399894
rect 278234 399574 278854 399658
rect 278234 399338 278266 399574
rect 278502 399338 278586 399574
rect 278822 399338 278854 399574
rect 278234 339894 278854 399338
rect 278234 339658 278266 339894
rect 278502 339658 278586 339894
rect 278822 339658 278854 339894
rect 278234 339574 278854 339658
rect 278234 339338 278266 339574
rect 278502 339338 278586 339574
rect 278822 339338 278854 339574
rect 278234 279894 278854 339338
rect 278234 279658 278266 279894
rect 278502 279658 278586 279894
rect 278822 279658 278854 279894
rect 278234 279574 278854 279658
rect 278234 279338 278266 279574
rect 278502 279338 278586 279574
rect 278822 279338 278854 279574
rect 278234 219894 278854 279338
rect 278234 219658 278266 219894
rect 278502 219658 278586 219894
rect 278822 219658 278854 219894
rect 278234 219574 278854 219658
rect 278234 219338 278266 219574
rect 278502 219338 278586 219574
rect 278822 219338 278854 219574
rect 278234 159894 278854 219338
rect 278234 159658 278266 159894
rect 278502 159658 278586 159894
rect 278822 159658 278854 159894
rect 278234 159574 278854 159658
rect 278234 159338 278266 159574
rect 278502 159338 278586 159574
rect 278822 159338 278854 159574
rect 278234 99894 278854 159338
rect 278234 99658 278266 99894
rect 278502 99658 278586 99894
rect 278822 99658 278854 99894
rect 278234 99574 278854 99658
rect 278234 99338 278266 99574
rect 278502 99338 278586 99574
rect 278822 99338 278854 99574
rect 278234 39894 278854 99338
rect 278234 39658 278266 39894
rect 278502 39658 278586 39894
rect 278822 39658 278854 39894
rect 278234 39574 278854 39658
rect 278234 39338 278266 39574
rect 278502 39338 278586 39574
rect 278822 39338 278854 39574
rect 278234 -5146 278854 39338
rect 278234 -5382 278266 -5146
rect 278502 -5382 278586 -5146
rect 278822 -5382 278854 -5146
rect 278234 -5466 278854 -5382
rect 278234 -5702 278266 -5466
rect 278502 -5702 278586 -5466
rect 278822 -5702 278854 -5466
rect 278234 -5734 278854 -5702
rect 281954 643614 282574 711002
rect 311954 710598 312574 711590
rect 311954 710362 311986 710598
rect 312222 710362 312306 710598
rect 312542 710362 312574 710598
rect 311954 710278 312574 710362
rect 311954 710042 311986 710278
rect 312222 710042 312306 710278
rect 312542 710042 312574 710278
rect 308234 708678 308854 709670
rect 308234 708442 308266 708678
rect 308502 708442 308586 708678
rect 308822 708442 308854 708678
rect 308234 708358 308854 708442
rect 308234 708122 308266 708358
rect 308502 708122 308586 708358
rect 308822 708122 308854 708358
rect 304514 706758 305134 707750
rect 304514 706522 304546 706758
rect 304782 706522 304866 706758
rect 305102 706522 305134 706758
rect 304514 706438 305134 706522
rect 304514 706202 304546 706438
rect 304782 706202 304866 706438
rect 305102 706202 305134 706438
rect 281954 643378 281986 643614
rect 282222 643378 282306 643614
rect 282542 643378 282574 643614
rect 281954 643294 282574 643378
rect 281954 643058 281986 643294
rect 282222 643058 282306 643294
rect 282542 643058 282574 643294
rect 281954 583614 282574 643058
rect 281954 583378 281986 583614
rect 282222 583378 282306 583614
rect 282542 583378 282574 583614
rect 281954 583294 282574 583378
rect 281954 583058 281986 583294
rect 282222 583058 282306 583294
rect 282542 583058 282574 583294
rect 281954 523614 282574 583058
rect 281954 523378 281986 523614
rect 282222 523378 282306 523614
rect 282542 523378 282574 523614
rect 281954 523294 282574 523378
rect 281954 523058 281986 523294
rect 282222 523058 282306 523294
rect 282542 523058 282574 523294
rect 281954 463614 282574 523058
rect 281954 463378 281986 463614
rect 282222 463378 282306 463614
rect 282542 463378 282574 463614
rect 281954 463294 282574 463378
rect 281954 463058 281986 463294
rect 282222 463058 282306 463294
rect 282542 463058 282574 463294
rect 281954 403614 282574 463058
rect 281954 403378 281986 403614
rect 282222 403378 282306 403614
rect 282542 403378 282574 403614
rect 281954 403294 282574 403378
rect 281954 403058 281986 403294
rect 282222 403058 282306 403294
rect 282542 403058 282574 403294
rect 281954 343614 282574 403058
rect 281954 343378 281986 343614
rect 282222 343378 282306 343614
rect 282542 343378 282574 343614
rect 281954 343294 282574 343378
rect 281954 343058 281986 343294
rect 282222 343058 282306 343294
rect 282542 343058 282574 343294
rect 281954 283614 282574 343058
rect 281954 283378 281986 283614
rect 282222 283378 282306 283614
rect 282542 283378 282574 283614
rect 281954 283294 282574 283378
rect 281954 283058 281986 283294
rect 282222 283058 282306 283294
rect 282542 283058 282574 283294
rect 281954 223614 282574 283058
rect 281954 223378 281986 223614
rect 282222 223378 282306 223614
rect 282542 223378 282574 223614
rect 281954 223294 282574 223378
rect 281954 223058 281986 223294
rect 282222 223058 282306 223294
rect 282542 223058 282574 223294
rect 281954 163614 282574 223058
rect 281954 163378 281986 163614
rect 282222 163378 282306 163614
rect 282542 163378 282574 163614
rect 281954 163294 282574 163378
rect 281954 163058 281986 163294
rect 282222 163058 282306 163294
rect 282542 163058 282574 163294
rect 281954 103614 282574 163058
rect 281954 103378 281986 103614
rect 282222 103378 282306 103614
rect 282542 103378 282574 103614
rect 281954 103294 282574 103378
rect 281954 103058 281986 103294
rect 282222 103058 282306 103294
rect 282542 103058 282574 103294
rect 281954 43614 282574 103058
rect 281954 43378 281986 43614
rect 282222 43378 282306 43614
rect 282542 43378 282574 43614
rect 281954 43294 282574 43378
rect 281954 43058 281986 43294
rect 282222 43058 282306 43294
rect 282542 43058 282574 43294
rect 251954 -6342 251986 -6106
rect 252222 -6342 252306 -6106
rect 252542 -6342 252574 -6106
rect 251954 -6426 252574 -6342
rect 251954 -6662 251986 -6426
rect 252222 -6662 252306 -6426
rect 252542 -6662 252574 -6426
rect 251954 -7654 252574 -6662
rect 281954 -7066 282574 43058
rect 300794 704838 301414 705830
rect 300794 704602 300826 704838
rect 301062 704602 301146 704838
rect 301382 704602 301414 704838
rect 300794 704518 301414 704602
rect 300794 704282 300826 704518
rect 301062 704282 301146 704518
rect 301382 704282 301414 704518
rect 300794 662454 301414 704282
rect 300794 662218 300826 662454
rect 301062 662218 301146 662454
rect 301382 662218 301414 662454
rect 300794 662134 301414 662218
rect 300794 661898 300826 662134
rect 301062 661898 301146 662134
rect 301382 661898 301414 662134
rect 300794 602454 301414 661898
rect 300794 602218 300826 602454
rect 301062 602218 301146 602454
rect 301382 602218 301414 602454
rect 300794 602134 301414 602218
rect 300794 601898 300826 602134
rect 301062 601898 301146 602134
rect 301382 601898 301414 602134
rect 300794 542454 301414 601898
rect 300794 542218 300826 542454
rect 301062 542218 301146 542454
rect 301382 542218 301414 542454
rect 300794 542134 301414 542218
rect 300794 541898 300826 542134
rect 301062 541898 301146 542134
rect 301382 541898 301414 542134
rect 300794 482454 301414 541898
rect 300794 482218 300826 482454
rect 301062 482218 301146 482454
rect 301382 482218 301414 482454
rect 300794 482134 301414 482218
rect 300794 481898 300826 482134
rect 301062 481898 301146 482134
rect 301382 481898 301414 482134
rect 300794 422454 301414 481898
rect 300794 422218 300826 422454
rect 301062 422218 301146 422454
rect 301382 422218 301414 422454
rect 300794 422134 301414 422218
rect 300794 421898 300826 422134
rect 301062 421898 301146 422134
rect 301382 421898 301414 422134
rect 300794 362454 301414 421898
rect 300794 362218 300826 362454
rect 301062 362218 301146 362454
rect 301382 362218 301414 362454
rect 300794 362134 301414 362218
rect 300794 361898 300826 362134
rect 301062 361898 301146 362134
rect 301382 361898 301414 362134
rect 300794 302454 301414 361898
rect 300794 302218 300826 302454
rect 301062 302218 301146 302454
rect 301382 302218 301414 302454
rect 300794 302134 301414 302218
rect 300794 301898 300826 302134
rect 301062 301898 301146 302134
rect 301382 301898 301414 302134
rect 300794 242454 301414 301898
rect 300794 242218 300826 242454
rect 301062 242218 301146 242454
rect 301382 242218 301414 242454
rect 300794 242134 301414 242218
rect 300794 241898 300826 242134
rect 301062 241898 301146 242134
rect 301382 241898 301414 242134
rect 300794 182454 301414 241898
rect 300794 182218 300826 182454
rect 301062 182218 301146 182454
rect 301382 182218 301414 182454
rect 300794 182134 301414 182218
rect 300794 181898 300826 182134
rect 301062 181898 301146 182134
rect 301382 181898 301414 182134
rect 300794 122454 301414 181898
rect 300794 122218 300826 122454
rect 301062 122218 301146 122454
rect 301382 122218 301414 122454
rect 300794 122134 301414 122218
rect 300794 121898 300826 122134
rect 301062 121898 301146 122134
rect 301382 121898 301414 122134
rect 300794 62454 301414 121898
rect 300794 62218 300826 62454
rect 301062 62218 301146 62454
rect 301382 62218 301414 62454
rect 300794 62134 301414 62218
rect 300794 61898 300826 62134
rect 301062 61898 301146 62134
rect 301382 61898 301414 62134
rect 300794 2454 301414 61898
rect 300794 2218 300826 2454
rect 301062 2218 301146 2454
rect 301382 2218 301414 2454
rect 300794 2134 301414 2218
rect 300794 1898 300826 2134
rect 301062 1898 301146 2134
rect 301382 1898 301414 2134
rect 300794 -346 301414 1898
rect 300794 -582 300826 -346
rect 301062 -582 301146 -346
rect 301382 -582 301414 -346
rect 300794 -666 301414 -582
rect 300794 -902 300826 -666
rect 301062 -902 301146 -666
rect 301382 -902 301414 -666
rect 300794 -1894 301414 -902
rect 304514 666174 305134 706202
rect 304514 665938 304546 666174
rect 304782 665938 304866 666174
rect 305102 665938 305134 666174
rect 304514 665854 305134 665938
rect 304514 665618 304546 665854
rect 304782 665618 304866 665854
rect 305102 665618 305134 665854
rect 304514 606174 305134 665618
rect 304514 605938 304546 606174
rect 304782 605938 304866 606174
rect 305102 605938 305134 606174
rect 304514 605854 305134 605938
rect 304514 605618 304546 605854
rect 304782 605618 304866 605854
rect 305102 605618 305134 605854
rect 304514 546174 305134 605618
rect 304514 545938 304546 546174
rect 304782 545938 304866 546174
rect 305102 545938 305134 546174
rect 304514 545854 305134 545938
rect 304514 545618 304546 545854
rect 304782 545618 304866 545854
rect 305102 545618 305134 545854
rect 304514 486174 305134 545618
rect 304514 485938 304546 486174
rect 304782 485938 304866 486174
rect 305102 485938 305134 486174
rect 304514 485854 305134 485938
rect 304514 485618 304546 485854
rect 304782 485618 304866 485854
rect 305102 485618 305134 485854
rect 304514 426174 305134 485618
rect 304514 425938 304546 426174
rect 304782 425938 304866 426174
rect 305102 425938 305134 426174
rect 304514 425854 305134 425938
rect 304514 425618 304546 425854
rect 304782 425618 304866 425854
rect 305102 425618 305134 425854
rect 304514 366174 305134 425618
rect 304514 365938 304546 366174
rect 304782 365938 304866 366174
rect 305102 365938 305134 366174
rect 304514 365854 305134 365938
rect 304514 365618 304546 365854
rect 304782 365618 304866 365854
rect 305102 365618 305134 365854
rect 304514 306174 305134 365618
rect 304514 305938 304546 306174
rect 304782 305938 304866 306174
rect 305102 305938 305134 306174
rect 304514 305854 305134 305938
rect 304514 305618 304546 305854
rect 304782 305618 304866 305854
rect 305102 305618 305134 305854
rect 304514 246174 305134 305618
rect 304514 245938 304546 246174
rect 304782 245938 304866 246174
rect 305102 245938 305134 246174
rect 304514 245854 305134 245938
rect 304514 245618 304546 245854
rect 304782 245618 304866 245854
rect 305102 245618 305134 245854
rect 304514 186174 305134 245618
rect 304514 185938 304546 186174
rect 304782 185938 304866 186174
rect 305102 185938 305134 186174
rect 304514 185854 305134 185938
rect 304514 185618 304546 185854
rect 304782 185618 304866 185854
rect 305102 185618 305134 185854
rect 304514 126174 305134 185618
rect 304514 125938 304546 126174
rect 304782 125938 304866 126174
rect 305102 125938 305134 126174
rect 304514 125854 305134 125938
rect 304514 125618 304546 125854
rect 304782 125618 304866 125854
rect 305102 125618 305134 125854
rect 304514 66174 305134 125618
rect 304514 65938 304546 66174
rect 304782 65938 304866 66174
rect 305102 65938 305134 66174
rect 304514 65854 305134 65938
rect 304514 65618 304546 65854
rect 304782 65618 304866 65854
rect 305102 65618 305134 65854
rect 304514 6174 305134 65618
rect 304514 5938 304546 6174
rect 304782 5938 304866 6174
rect 305102 5938 305134 6174
rect 304514 5854 305134 5938
rect 304514 5618 304546 5854
rect 304782 5618 304866 5854
rect 305102 5618 305134 5854
rect 304514 -2266 305134 5618
rect 304514 -2502 304546 -2266
rect 304782 -2502 304866 -2266
rect 305102 -2502 305134 -2266
rect 304514 -2586 305134 -2502
rect 304514 -2822 304546 -2586
rect 304782 -2822 304866 -2586
rect 305102 -2822 305134 -2586
rect 304514 -3814 305134 -2822
rect 308234 669894 308854 708122
rect 308234 669658 308266 669894
rect 308502 669658 308586 669894
rect 308822 669658 308854 669894
rect 308234 669574 308854 669658
rect 308234 669338 308266 669574
rect 308502 669338 308586 669574
rect 308822 669338 308854 669574
rect 308234 609894 308854 669338
rect 308234 609658 308266 609894
rect 308502 609658 308586 609894
rect 308822 609658 308854 609894
rect 308234 609574 308854 609658
rect 308234 609338 308266 609574
rect 308502 609338 308586 609574
rect 308822 609338 308854 609574
rect 308234 549894 308854 609338
rect 308234 549658 308266 549894
rect 308502 549658 308586 549894
rect 308822 549658 308854 549894
rect 308234 549574 308854 549658
rect 308234 549338 308266 549574
rect 308502 549338 308586 549574
rect 308822 549338 308854 549574
rect 308234 489894 308854 549338
rect 308234 489658 308266 489894
rect 308502 489658 308586 489894
rect 308822 489658 308854 489894
rect 308234 489574 308854 489658
rect 308234 489338 308266 489574
rect 308502 489338 308586 489574
rect 308822 489338 308854 489574
rect 308234 429894 308854 489338
rect 308234 429658 308266 429894
rect 308502 429658 308586 429894
rect 308822 429658 308854 429894
rect 308234 429574 308854 429658
rect 308234 429338 308266 429574
rect 308502 429338 308586 429574
rect 308822 429338 308854 429574
rect 308234 369894 308854 429338
rect 308234 369658 308266 369894
rect 308502 369658 308586 369894
rect 308822 369658 308854 369894
rect 308234 369574 308854 369658
rect 308234 369338 308266 369574
rect 308502 369338 308586 369574
rect 308822 369338 308854 369574
rect 308234 309894 308854 369338
rect 308234 309658 308266 309894
rect 308502 309658 308586 309894
rect 308822 309658 308854 309894
rect 308234 309574 308854 309658
rect 308234 309338 308266 309574
rect 308502 309338 308586 309574
rect 308822 309338 308854 309574
rect 308234 249894 308854 309338
rect 308234 249658 308266 249894
rect 308502 249658 308586 249894
rect 308822 249658 308854 249894
rect 308234 249574 308854 249658
rect 308234 249338 308266 249574
rect 308502 249338 308586 249574
rect 308822 249338 308854 249574
rect 308234 189894 308854 249338
rect 308234 189658 308266 189894
rect 308502 189658 308586 189894
rect 308822 189658 308854 189894
rect 308234 189574 308854 189658
rect 308234 189338 308266 189574
rect 308502 189338 308586 189574
rect 308822 189338 308854 189574
rect 308234 129894 308854 189338
rect 308234 129658 308266 129894
rect 308502 129658 308586 129894
rect 308822 129658 308854 129894
rect 308234 129574 308854 129658
rect 308234 129338 308266 129574
rect 308502 129338 308586 129574
rect 308822 129338 308854 129574
rect 308234 69894 308854 129338
rect 308234 69658 308266 69894
rect 308502 69658 308586 69894
rect 308822 69658 308854 69894
rect 308234 69574 308854 69658
rect 308234 69338 308266 69574
rect 308502 69338 308586 69574
rect 308822 69338 308854 69574
rect 308234 9894 308854 69338
rect 308234 9658 308266 9894
rect 308502 9658 308586 9894
rect 308822 9658 308854 9894
rect 308234 9574 308854 9658
rect 308234 9338 308266 9574
rect 308502 9338 308586 9574
rect 308822 9338 308854 9574
rect 308234 -4186 308854 9338
rect 308234 -4422 308266 -4186
rect 308502 -4422 308586 -4186
rect 308822 -4422 308854 -4186
rect 308234 -4506 308854 -4422
rect 308234 -4742 308266 -4506
rect 308502 -4742 308586 -4506
rect 308822 -4742 308854 -4506
rect 308234 -5734 308854 -4742
rect 311954 673614 312574 710042
rect 341954 711558 342574 711590
rect 341954 711322 341986 711558
rect 342222 711322 342306 711558
rect 342542 711322 342574 711558
rect 341954 711238 342574 711322
rect 341954 711002 341986 711238
rect 342222 711002 342306 711238
rect 342542 711002 342574 711238
rect 338234 709638 338854 709670
rect 338234 709402 338266 709638
rect 338502 709402 338586 709638
rect 338822 709402 338854 709638
rect 338234 709318 338854 709402
rect 338234 709082 338266 709318
rect 338502 709082 338586 709318
rect 338822 709082 338854 709318
rect 334514 707718 335134 707750
rect 334514 707482 334546 707718
rect 334782 707482 334866 707718
rect 335102 707482 335134 707718
rect 334514 707398 335134 707482
rect 334514 707162 334546 707398
rect 334782 707162 334866 707398
rect 335102 707162 335134 707398
rect 311954 673378 311986 673614
rect 312222 673378 312306 673614
rect 312542 673378 312574 673614
rect 311954 673294 312574 673378
rect 311954 673058 311986 673294
rect 312222 673058 312306 673294
rect 312542 673058 312574 673294
rect 311954 613614 312574 673058
rect 311954 613378 311986 613614
rect 312222 613378 312306 613614
rect 312542 613378 312574 613614
rect 311954 613294 312574 613378
rect 311954 613058 311986 613294
rect 312222 613058 312306 613294
rect 312542 613058 312574 613294
rect 311954 553614 312574 613058
rect 311954 553378 311986 553614
rect 312222 553378 312306 553614
rect 312542 553378 312574 553614
rect 311954 553294 312574 553378
rect 311954 553058 311986 553294
rect 312222 553058 312306 553294
rect 312542 553058 312574 553294
rect 311954 493614 312574 553058
rect 311954 493378 311986 493614
rect 312222 493378 312306 493614
rect 312542 493378 312574 493614
rect 311954 493294 312574 493378
rect 311954 493058 311986 493294
rect 312222 493058 312306 493294
rect 312542 493058 312574 493294
rect 311954 433614 312574 493058
rect 311954 433378 311986 433614
rect 312222 433378 312306 433614
rect 312542 433378 312574 433614
rect 311954 433294 312574 433378
rect 311954 433058 311986 433294
rect 312222 433058 312306 433294
rect 312542 433058 312574 433294
rect 311954 373614 312574 433058
rect 311954 373378 311986 373614
rect 312222 373378 312306 373614
rect 312542 373378 312574 373614
rect 311954 373294 312574 373378
rect 311954 373058 311986 373294
rect 312222 373058 312306 373294
rect 312542 373058 312574 373294
rect 311954 313614 312574 373058
rect 311954 313378 311986 313614
rect 312222 313378 312306 313614
rect 312542 313378 312574 313614
rect 311954 313294 312574 313378
rect 311954 313058 311986 313294
rect 312222 313058 312306 313294
rect 312542 313058 312574 313294
rect 311954 253614 312574 313058
rect 311954 253378 311986 253614
rect 312222 253378 312306 253614
rect 312542 253378 312574 253614
rect 311954 253294 312574 253378
rect 311954 253058 311986 253294
rect 312222 253058 312306 253294
rect 312542 253058 312574 253294
rect 311954 193614 312574 253058
rect 311954 193378 311986 193614
rect 312222 193378 312306 193614
rect 312542 193378 312574 193614
rect 311954 193294 312574 193378
rect 311954 193058 311986 193294
rect 312222 193058 312306 193294
rect 312542 193058 312574 193294
rect 311954 133614 312574 193058
rect 311954 133378 311986 133614
rect 312222 133378 312306 133614
rect 312542 133378 312574 133614
rect 311954 133294 312574 133378
rect 311954 133058 311986 133294
rect 312222 133058 312306 133294
rect 312542 133058 312574 133294
rect 311954 73614 312574 133058
rect 311954 73378 311986 73614
rect 312222 73378 312306 73614
rect 312542 73378 312574 73614
rect 311954 73294 312574 73378
rect 311954 73058 311986 73294
rect 312222 73058 312306 73294
rect 312542 73058 312574 73294
rect 311954 13614 312574 73058
rect 311954 13378 311986 13614
rect 312222 13378 312306 13614
rect 312542 13378 312574 13614
rect 311954 13294 312574 13378
rect 311954 13058 311986 13294
rect 312222 13058 312306 13294
rect 312542 13058 312574 13294
rect 281954 -7302 281986 -7066
rect 282222 -7302 282306 -7066
rect 282542 -7302 282574 -7066
rect 281954 -7386 282574 -7302
rect 281954 -7622 281986 -7386
rect 282222 -7622 282306 -7386
rect 282542 -7622 282574 -7386
rect 281954 -7654 282574 -7622
rect 311954 -6106 312574 13058
rect 330794 705798 331414 705830
rect 330794 705562 330826 705798
rect 331062 705562 331146 705798
rect 331382 705562 331414 705798
rect 330794 705478 331414 705562
rect 330794 705242 330826 705478
rect 331062 705242 331146 705478
rect 331382 705242 331414 705478
rect 330794 692454 331414 705242
rect 330794 692218 330826 692454
rect 331062 692218 331146 692454
rect 331382 692218 331414 692454
rect 330794 692134 331414 692218
rect 330794 691898 330826 692134
rect 331062 691898 331146 692134
rect 331382 691898 331414 692134
rect 330794 632454 331414 691898
rect 330794 632218 330826 632454
rect 331062 632218 331146 632454
rect 331382 632218 331414 632454
rect 330794 632134 331414 632218
rect 330794 631898 330826 632134
rect 331062 631898 331146 632134
rect 331382 631898 331414 632134
rect 330794 572454 331414 631898
rect 330794 572218 330826 572454
rect 331062 572218 331146 572454
rect 331382 572218 331414 572454
rect 330794 572134 331414 572218
rect 330794 571898 330826 572134
rect 331062 571898 331146 572134
rect 331382 571898 331414 572134
rect 330794 512454 331414 571898
rect 330794 512218 330826 512454
rect 331062 512218 331146 512454
rect 331382 512218 331414 512454
rect 330794 512134 331414 512218
rect 330794 511898 330826 512134
rect 331062 511898 331146 512134
rect 331382 511898 331414 512134
rect 330794 452454 331414 511898
rect 330794 452218 330826 452454
rect 331062 452218 331146 452454
rect 331382 452218 331414 452454
rect 330794 452134 331414 452218
rect 330794 451898 330826 452134
rect 331062 451898 331146 452134
rect 331382 451898 331414 452134
rect 330794 392454 331414 451898
rect 330794 392218 330826 392454
rect 331062 392218 331146 392454
rect 331382 392218 331414 392454
rect 330794 392134 331414 392218
rect 330794 391898 330826 392134
rect 331062 391898 331146 392134
rect 331382 391898 331414 392134
rect 330794 332454 331414 391898
rect 330794 332218 330826 332454
rect 331062 332218 331146 332454
rect 331382 332218 331414 332454
rect 330794 332134 331414 332218
rect 330794 331898 330826 332134
rect 331062 331898 331146 332134
rect 331382 331898 331414 332134
rect 330794 272454 331414 331898
rect 330794 272218 330826 272454
rect 331062 272218 331146 272454
rect 331382 272218 331414 272454
rect 330794 272134 331414 272218
rect 330794 271898 330826 272134
rect 331062 271898 331146 272134
rect 331382 271898 331414 272134
rect 330794 212454 331414 271898
rect 330794 212218 330826 212454
rect 331062 212218 331146 212454
rect 331382 212218 331414 212454
rect 330794 212134 331414 212218
rect 330794 211898 330826 212134
rect 331062 211898 331146 212134
rect 331382 211898 331414 212134
rect 330794 152454 331414 211898
rect 330794 152218 330826 152454
rect 331062 152218 331146 152454
rect 331382 152218 331414 152454
rect 330794 152134 331414 152218
rect 330794 151898 330826 152134
rect 331062 151898 331146 152134
rect 331382 151898 331414 152134
rect 330794 92454 331414 151898
rect 330794 92218 330826 92454
rect 331062 92218 331146 92454
rect 331382 92218 331414 92454
rect 330794 92134 331414 92218
rect 330794 91898 330826 92134
rect 331062 91898 331146 92134
rect 331382 91898 331414 92134
rect 330794 32454 331414 91898
rect 330794 32218 330826 32454
rect 331062 32218 331146 32454
rect 331382 32218 331414 32454
rect 330794 32134 331414 32218
rect 330794 31898 330826 32134
rect 331062 31898 331146 32134
rect 331382 31898 331414 32134
rect 330794 -1306 331414 31898
rect 330794 -1542 330826 -1306
rect 331062 -1542 331146 -1306
rect 331382 -1542 331414 -1306
rect 330794 -1626 331414 -1542
rect 330794 -1862 330826 -1626
rect 331062 -1862 331146 -1626
rect 331382 -1862 331414 -1626
rect 330794 -1894 331414 -1862
rect 334514 696174 335134 707162
rect 334514 695938 334546 696174
rect 334782 695938 334866 696174
rect 335102 695938 335134 696174
rect 334514 695854 335134 695938
rect 334514 695618 334546 695854
rect 334782 695618 334866 695854
rect 335102 695618 335134 695854
rect 334514 636174 335134 695618
rect 334514 635938 334546 636174
rect 334782 635938 334866 636174
rect 335102 635938 335134 636174
rect 334514 635854 335134 635938
rect 334514 635618 334546 635854
rect 334782 635618 334866 635854
rect 335102 635618 335134 635854
rect 334514 576174 335134 635618
rect 334514 575938 334546 576174
rect 334782 575938 334866 576174
rect 335102 575938 335134 576174
rect 334514 575854 335134 575938
rect 334514 575618 334546 575854
rect 334782 575618 334866 575854
rect 335102 575618 335134 575854
rect 334514 516174 335134 575618
rect 334514 515938 334546 516174
rect 334782 515938 334866 516174
rect 335102 515938 335134 516174
rect 334514 515854 335134 515938
rect 334514 515618 334546 515854
rect 334782 515618 334866 515854
rect 335102 515618 335134 515854
rect 334514 456174 335134 515618
rect 334514 455938 334546 456174
rect 334782 455938 334866 456174
rect 335102 455938 335134 456174
rect 334514 455854 335134 455938
rect 334514 455618 334546 455854
rect 334782 455618 334866 455854
rect 335102 455618 335134 455854
rect 334514 396174 335134 455618
rect 334514 395938 334546 396174
rect 334782 395938 334866 396174
rect 335102 395938 335134 396174
rect 334514 395854 335134 395938
rect 334514 395618 334546 395854
rect 334782 395618 334866 395854
rect 335102 395618 335134 395854
rect 334514 336174 335134 395618
rect 334514 335938 334546 336174
rect 334782 335938 334866 336174
rect 335102 335938 335134 336174
rect 334514 335854 335134 335938
rect 334514 335618 334546 335854
rect 334782 335618 334866 335854
rect 335102 335618 335134 335854
rect 334514 276174 335134 335618
rect 334514 275938 334546 276174
rect 334782 275938 334866 276174
rect 335102 275938 335134 276174
rect 334514 275854 335134 275938
rect 334514 275618 334546 275854
rect 334782 275618 334866 275854
rect 335102 275618 335134 275854
rect 334514 216174 335134 275618
rect 334514 215938 334546 216174
rect 334782 215938 334866 216174
rect 335102 215938 335134 216174
rect 334514 215854 335134 215938
rect 334514 215618 334546 215854
rect 334782 215618 334866 215854
rect 335102 215618 335134 215854
rect 334514 156174 335134 215618
rect 334514 155938 334546 156174
rect 334782 155938 334866 156174
rect 335102 155938 335134 156174
rect 334514 155854 335134 155938
rect 334514 155618 334546 155854
rect 334782 155618 334866 155854
rect 335102 155618 335134 155854
rect 334514 96174 335134 155618
rect 334514 95938 334546 96174
rect 334782 95938 334866 96174
rect 335102 95938 335134 96174
rect 334514 95854 335134 95938
rect 334514 95618 334546 95854
rect 334782 95618 334866 95854
rect 335102 95618 335134 95854
rect 334514 36174 335134 95618
rect 334514 35938 334546 36174
rect 334782 35938 334866 36174
rect 335102 35938 335134 36174
rect 334514 35854 335134 35938
rect 334514 35618 334546 35854
rect 334782 35618 334866 35854
rect 335102 35618 335134 35854
rect 334514 -3226 335134 35618
rect 334514 -3462 334546 -3226
rect 334782 -3462 334866 -3226
rect 335102 -3462 335134 -3226
rect 334514 -3546 335134 -3462
rect 334514 -3782 334546 -3546
rect 334782 -3782 334866 -3546
rect 335102 -3782 335134 -3546
rect 334514 -3814 335134 -3782
rect 338234 699894 338854 709082
rect 338234 699658 338266 699894
rect 338502 699658 338586 699894
rect 338822 699658 338854 699894
rect 338234 699574 338854 699658
rect 338234 699338 338266 699574
rect 338502 699338 338586 699574
rect 338822 699338 338854 699574
rect 338234 639894 338854 699338
rect 338234 639658 338266 639894
rect 338502 639658 338586 639894
rect 338822 639658 338854 639894
rect 338234 639574 338854 639658
rect 338234 639338 338266 639574
rect 338502 639338 338586 639574
rect 338822 639338 338854 639574
rect 338234 579894 338854 639338
rect 338234 579658 338266 579894
rect 338502 579658 338586 579894
rect 338822 579658 338854 579894
rect 338234 579574 338854 579658
rect 338234 579338 338266 579574
rect 338502 579338 338586 579574
rect 338822 579338 338854 579574
rect 338234 519894 338854 579338
rect 338234 519658 338266 519894
rect 338502 519658 338586 519894
rect 338822 519658 338854 519894
rect 338234 519574 338854 519658
rect 338234 519338 338266 519574
rect 338502 519338 338586 519574
rect 338822 519338 338854 519574
rect 338234 459894 338854 519338
rect 338234 459658 338266 459894
rect 338502 459658 338586 459894
rect 338822 459658 338854 459894
rect 338234 459574 338854 459658
rect 338234 459338 338266 459574
rect 338502 459338 338586 459574
rect 338822 459338 338854 459574
rect 338234 399894 338854 459338
rect 338234 399658 338266 399894
rect 338502 399658 338586 399894
rect 338822 399658 338854 399894
rect 338234 399574 338854 399658
rect 338234 399338 338266 399574
rect 338502 399338 338586 399574
rect 338822 399338 338854 399574
rect 338234 339894 338854 399338
rect 338234 339658 338266 339894
rect 338502 339658 338586 339894
rect 338822 339658 338854 339894
rect 338234 339574 338854 339658
rect 338234 339338 338266 339574
rect 338502 339338 338586 339574
rect 338822 339338 338854 339574
rect 338234 279894 338854 339338
rect 338234 279658 338266 279894
rect 338502 279658 338586 279894
rect 338822 279658 338854 279894
rect 338234 279574 338854 279658
rect 338234 279338 338266 279574
rect 338502 279338 338586 279574
rect 338822 279338 338854 279574
rect 338234 219894 338854 279338
rect 338234 219658 338266 219894
rect 338502 219658 338586 219894
rect 338822 219658 338854 219894
rect 338234 219574 338854 219658
rect 338234 219338 338266 219574
rect 338502 219338 338586 219574
rect 338822 219338 338854 219574
rect 338234 159894 338854 219338
rect 338234 159658 338266 159894
rect 338502 159658 338586 159894
rect 338822 159658 338854 159894
rect 338234 159574 338854 159658
rect 338234 159338 338266 159574
rect 338502 159338 338586 159574
rect 338822 159338 338854 159574
rect 338234 99894 338854 159338
rect 338234 99658 338266 99894
rect 338502 99658 338586 99894
rect 338822 99658 338854 99894
rect 338234 99574 338854 99658
rect 338234 99338 338266 99574
rect 338502 99338 338586 99574
rect 338822 99338 338854 99574
rect 338234 39894 338854 99338
rect 338234 39658 338266 39894
rect 338502 39658 338586 39894
rect 338822 39658 338854 39894
rect 338234 39574 338854 39658
rect 338234 39338 338266 39574
rect 338502 39338 338586 39574
rect 338822 39338 338854 39574
rect 338234 -5146 338854 39338
rect 338234 -5382 338266 -5146
rect 338502 -5382 338586 -5146
rect 338822 -5382 338854 -5146
rect 338234 -5466 338854 -5382
rect 338234 -5702 338266 -5466
rect 338502 -5702 338586 -5466
rect 338822 -5702 338854 -5466
rect 338234 -5734 338854 -5702
rect 341954 643614 342574 711002
rect 371954 710598 372574 711590
rect 371954 710362 371986 710598
rect 372222 710362 372306 710598
rect 372542 710362 372574 710598
rect 371954 710278 372574 710362
rect 371954 710042 371986 710278
rect 372222 710042 372306 710278
rect 372542 710042 372574 710278
rect 368234 708678 368854 709670
rect 368234 708442 368266 708678
rect 368502 708442 368586 708678
rect 368822 708442 368854 708678
rect 368234 708358 368854 708442
rect 368234 708122 368266 708358
rect 368502 708122 368586 708358
rect 368822 708122 368854 708358
rect 364514 706758 365134 707750
rect 364514 706522 364546 706758
rect 364782 706522 364866 706758
rect 365102 706522 365134 706758
rect 364514 706438 365134 706522
rect 364514 706202 364546 706438
rect 364782 706202 364866 706438
rect 365102 706202 365134 706438
rect 341954 643378 341986 643614
rect 342222 643378 342306 643614
rect 342542 643378 342574 643614
rect 341954 643294 342574 643378
rect 341954 643058 341986 643294
rect 342222 643058 342306 643294
rect 342542 643058 342574 643294
rect 341954 583614 342574 643058
rect 341954 583378 341986 583614
rect 342222 583378 342306 583614
rect 342542 583378 342574 583614
rect 341954 583294 342574 583378
rect 341954 583058 341986 583294
rect 342222 583058 342306 583294
rect 342542 583058 342574 583294
rect 341954 523614 342574 583058
rect 341954 523378 341986 523614
rect 342222 523378 342306 523614
rect 342542 523378 342574 523614
rect 341954 523294 342574 523378
rect 341954 523058 341986 523294
rect 342222 523058 342306 523294
rect 342542 523058 342574 523294
rect 341954 463614 342574 523058
rect 341954 463378 341986 463614
rect 342222 463378 342306 463614
rect 342542 463378 342574 463614
rect 341954 463294 342574 463378
rect 341954 463058 341986 463294
rect 342222 463058 342306 463294
rect 342542 463058 342574 463294
rect 341954 403614 342574 463058
rect 341954 403378 341986 403614
rect 342222 403378 342306 403614
rect 342542 403378 342574 403614
rect 341954 403294 342574 403378
rect 341954 403058 341986 403294
rect 342222 403058 342306 403294
rect 342542 403058 342574 403294
rect 341954 343614 342574 403058
rect 341954 343378 341986 343614
rect 342222 343378 342306 343614
rect 342542 343378 342574 343614
rect 341954 343294 342574 343378
rect 341954 343058 341986 343294
rect 342222 343058 342306 343294
rect 342542 343058 342574 343294
rect 341954 283614 342574 343058
rect 341954 283378 341986 283614
rect 342222 283378 342306 283614
rect 342542 283378 342574 283614
rect 341954 283294 342574 283378
rect 341954 283058 341986 283294
rect 342222 283058 342306 283294
rect 342542 283058 342574 283294
rect 341954 223614 342574 283058
rect 341954 223378 341986 223614
rect 342222 223378 342306 223614
rect 342542 223378 342574 223614
rect 341954 223294 342574 223378
rect 341954 223058 341986 223294
rect 342222 223058 342306 223294
rect 342542 223058 342574 223294
rect 341954 163614 342574 223058
rect 341954 163378 341986 163614
rect 342222 163378 342306 163614
rect 342542 163378 342574 163614
rect 341954 163294 342574 163378
rect 341954 163058 341986 163294
rect 342222 163058 342306 163294
rect 342542 163058 342574 163294
rect 341954 103614 342574 163058
rect 341954 103378 341986 103614
rect 342222 103378 342306 103614
rect 342542 103378 342574 103614
rect 341954 103294 342574 103378
rect 341954 103058 341986 103294
rect 342222 103058 342306 103294
rect 342542 103058 342574 103294
rect 341954 43614 342574 103058
rect 341954 43378 341986 43614
rect 342222 43378 342306 43614
rect 342542 43378 342574 43614
rect 341954 43294 342574 43378
rect 341954 43058 341986 43294
rect 342222 43058 342306 43294
rect 342542 43058 342574 43294
rect 311954 -6342 311986 -6106
rect 312222 -6342 312306 -6106
rect 312542 -6342 312574 -6106
rect 311954 -6426 312574 -6342
rect 311954 -6662 311986 -6426
rect 312222 -6662 312306 -6426
rect 312542 -6662 312574 -6426
rect 311954 -7654 312574 -6662
rect 341954 -7066 342574 43058
rect 360794 704838 361414 705830
rect 360794 704602 360826 704838
rect 361062 704602 361146 704838
rect 361382 704602 361414 704838
rect 360794 704518 361414 704602
rect 360794 704282 360826 704518
rect 361062 704282 361146 704518
rect 361382 704282 361414 704518
rect 360794 662454 361414 704282
rect 360794 662218 360826 662454
rect 361062 662218 361146 662454
rect 361382 662218 361414 662454
rect 360794 662134 361414 662218
rect 360794 661898 360826 662134
rect 361062 661898 361146 662134
rect 361382 661898 361414 662134
rect 360794 602454 361414 661898
rect 360794 602218 360826 602454
rect 361062 602218 361146 602454
rect 361382 602218 361414 602454
rect 360794 602134 361414 602218
rect 360794 601898 360826 602134
rect 361062 601898 361146 602134
rect 361382 601898 361414 602134
rect 360794 542454 361414 601898
rect 360794 542218 360826 542454
rect 361062 542218 361146 542454
rect 361382 542218 361414 542454
rect 360794 542134 361414 542218
rect 360794 541898 360826 542134
rect 361062 541898 361146 542134
rect 361382 541898 361414 542134
rect 360794 482454 361414 541898
rect 360794 482218 360826 482454
rect 361062 482218 361146 482454
rect 361382 482218 361414 482454
rect 360794 482134 361414 482218
rect 360794 481898 360826 482134
rect 361062 481898 361146 482134
rect 361382 481898 361414 482134
rect 360794 422454 361414 481898
rect 360794 422218 360826 422454
rect 361062 422218 361146 422454
rect 361382 422218 361414 422454
rect 360794 422134 361414 422218
rect 360794 421898 360826 422134
rect 361062 421898 361146 422134
rect 361382 421898 361414 422134
rect 360794 362454 361414 421898
rect 360794 362218 360826 362454
rect 361062 362218 361146 362454
rect 361382 362218 361414 362454
rect 360794 362134 361414 362218
rect 360794 361898 360826 362134
rect 361062 361898 361146 362134
rect 361382 361898 361414 362134
rect 360794 302454 361414 361898
rect 360794 302218 360826 302454
rect 361062 302218 361146 302454
rect 361382 302218 361414 302454
rect 360794 302134 361414 302218
rect 360794 301898 360826 302134
rect 361062 301898 361146 302134
rect 361382 301898 361414 302134
rect 360794 242454 361414 301898
rect 360794 242218 360826 242454
rect 361062 242218 361146 242454
rect 361382 242218 361414 242454
rect 360794 242134 361414 242218
rect 360794 241898 360826 242134
rect 361062 241898 361146 242134
rect 361382 241898 361414 242134
rect 360794 182454 361414 241898
rect 360794 182218 360826 182454
rect 361062 182218 361146 182454
rect 361382 182218 361414 182454
rect 360794 182134 361414 182218
rect 360794 181898 360826 182134
rect 361062 181898 361146 182134
rect 361382 181898 361414 182134
rect 360794 122454 361414 181898
rect 360794 122218 360826 122454
rect 361062 122218 361146 122454
rect 361382 122218 361414 122454
rect 360794 122134 361414 122218
rect 360794 121898 360826 122134
rect 361062 121898 361146 122134
rect 361382 121898 361414 122134
rect 360794 62454 361414 121898
rect 360794 62218 360826 62454
rect 361062 62218 361146 62454
rect 361382 62218 361414 62454
rect 360794 62134 361414 62218
rect 360794 61898 360826 62134
rect 361062 61898 361146 62134
rect 361382 61898 361414 62134
rect 360794 2454 361414 61898
rect 360794 2218 360826 2454
rect 361062 2218 361146 2454
rect 361382 2218 361414 2454
rect 360794 2134 361414 2218
rect 360794 1898 360826 2134
rect 361062 1898 361146 2134
rect 361382 1898 361414 2134
rect 360794 -346 361414 1898
rect 360794 -582 360826 -346
rect 361062 -582 361146 -346
rect 361382 -582 361414 -346
rect 360794 -666 361414 -582
rect 360794 -902 360826 -666
rect 361062 -902 361146 -666
rect 361382 -902 361414 -666
rect 360794 -1894 361414 -902
rect 364514 666174 365134 706202
rect 364514 665938 364546 666174
rect 364782 665938 364866 666174
rect 365102 665938 365134 666174
rect 364514 665854 365134 665938
rect 364514 665618 364546 665854
rect 364782 665618 364866 665854
rect 365102 665618 365134 665854
rect 364514 606174 365134 665618
rect 364514 605938 364546 606174
rect 364782 605938 364866 606174
rect 365102 605938 365134 606174
rect 364514 605854 365134 605938
rect 364514 605618 364546 605854
rect 364782 605618 364866 605854
rect 365102 605618 365134 605854
rect 364514 546174 365134 605618
rect 364514 545938 364546 546174
rect 364782 545938 364866 546174
rect 365102 545938 365134 546174
rect 364514 545854 365134 545938
rect 364514 545618 364546 545854
rect 364782 545618 364866 545854
rect 365102 545618 365134 545854
rect 364514 486174 365134 545618
rect 364514 485938 364546 486174
rect 364782 485938 364866 486174
rect 365102 485938 365134 486174
rect 364514 485854 365134 485938
rect 364514 485618 364546 485854
rect 364782 485618 364866 485854
rect 365102 485618 365134 485854
rect 364514 426174 365134 485618
rect 364514 425938 364546 426174
rect 364782 425938 364866 426174
rect 365102 425938 365134 426174
rect 364514 425854 365134 425938
rect 364514 425618 364546 425854
rect 364782 425618 364866 425854
rect 365102 425618 365134 425854
rect 364514 366174 365134 425618
rect 364514 365938 364546 366174
rect 364782 365938 364866 366174
rect 365102 365938 365134 366174
rect 364514 365854 365134 365938
rect 364514 365618 364546 365854
rect 364782 365618 364866 365854
rect 365102 365618 365134 365854
rect 364514 306174 365134 365618
rect 364514 305938 364546 306174
rect 364782 305938 364866 306174
rect 365102 305938 365134 306174
rect 364514 305854 365134 305938
rect 364514 305618 364546 305854
rect 364782 305618 364866 305854
rect 365102 305618 365134 305854
rect 364514 246174 365134 305618
rect 364514 245938 364546 246174
rect 364782 245938 364866 246174
rect 365102 245938 365134 246174
rect 364514 245854 365134 245938
rect 364514 245618 364546 245854
rect 364782 245618 364866 245854
rect 365102 245618 365134 245854
rect 364514 186174 365134 245618
rect 364514 185938 364546 186174
rect 364782 185938 364866 186174
rect 365102 185938 365134 186174
rect 364514 185854 365134 185938
rect 364514 185618 364546 185854
rect 364782 185618 364866 185854
rect 365102 185618 365134 185854
rect 364514 126174 365134 185618
rect 364514 125938 364546 126174
rect 364782 125938 364866 126174
rect 365102 125938 365134 126174
rect 364514 125854 365134 125938
rect 364514 125618 364546 125854
rect 364782 125618 364866 125854
rect 365102 125618 365134 125854
rect 364514 66174 365134 125618
rect 364514 65938 364546 66174
rect 364782 65938 364866 66174
rect 365102 65938 365134 66174
rect 364514 65854 365134 65938
rect 364514 65618 364546 65854
rect 364782 65618 364866 65854
rect 365102 65618 365134 65854
rect 364514 6174 365134 65618
rect 364514 5938 364546 6174
rect 364782 5938 364866 6174
rect 365102 5938 365134 6174
rect 364514 5854 365134 5938
rect 364514 5618 364546 5854
rect 364782 5618 364866 5854
rect 365102 5618 365134 5854
rect 364514 -2266 365134 5618
rect 364514 -2502 364546 -2266
rect 364782 -2502 364866 -2266
rect 365102 -2502 365134 -2266
rect 364514 -2586 365134 -2502
rect 364514 -2822 364546 -2586
rect 364782 -2822 364866 -2586
rect 365102 -2822 365134 -2586
rect 364514 -3814 365134 -2822
rect 368234 669894 368854 708122
rect 368234 669658 368266 669894
rect 368502 669658 368586 669894
rect 368822 669658 368854 669894
rect 368234 669574 368854 669658
rect 368234 669338 368266 669574
rect 368502 669338 368586 669574
rect 368822 669338 368854 669574
rect 368234 609894 368854 669338
rect 368234 609658 368266 609894
rect 368502 609658 368586 609894
rect 368822 609658 368854 609894
rect 368234 609574 368854 609658
rect 368234 609338 368266 609574
rect 368502 609338 368586 609574
rect 368822 609338 368854 609574
rect 368234 549894 368854 609338
rect 368234 549658 368266 549894
rect 368502 549658 368586 549894
rect 368822 549658 368854 549894
rect 368234 549574 368854 549658
rect 368234 549338 368266 549574
rect 368502 549338 368586 549574
rect 368822 549338 368854 549574
rect 368234 489894 368854 549338
rect 368234 489658 368266 489894
rect 368502 489658 368586 489894
rect 368822 489658 368854 489894
rect 368234 489574 368854 489658
rect 368234 489338 368266 489574
rect 368502 489338 368586 489574
rect 368822 489338 368854 489574
rect 368234 429894 368854 489338
rect 368234 429658 368266 429894
rect 368502 429658 368586 429894
rect 368822 429658 368854 429894
rect 368234 429574 368854 429658
rect 368234 429338 368266 429574
rect 368502 429338 368586 429574
rect 368822 429338 368854 429574
rect 368234 369894 368854 429338
rect 368234 369658 368266 369894
rect 368502 369658 368586 369894
rect 368822 369658 368854 369894
rect 368234 369574 368854 369658
rect 368234 369338 368266 369574
rect 368502 369338 368586 369574
rect 368822 369338 368854 369574
rect 368234 309894 368854 369338
rect 368234 309658 368266 309894
rect 368502 309658 368586 309894
rect 368822 309658 368854 309894
rect 368234 309574 368854 309658
rect 368234 309338 368266 309574
rect 368502 309338 368586 309574
rect 368822 309338 368854 309574
rect 368234 249894 368854 309338
rect 368234 249658 368266 249894
rect 368502 249658 368586 249894
rect 368822 249658 368854 249894
rect 368234 249574 368854 249658
rect 368234 249338 368266 249574
rect 368502 249338 368586 249574
rect 368822 249338 368854 249574
rect 368234 189894 368854 249338
rect 368234 189658 368266 189894
rect 368502 189658 368586 189894
rect 368822 189658 368854 189894
rect 368234 189574 368854 189658
rect 368234 189338 368266 189574
rect 368502 189338 368586 189574
rect 368822 189338 368854 189574
rect 368234 129894 368854 189338
rect 368234 129658 368266 129894
rect 368502 129658 368586 129894
rect 368822 129658 368854 129894
rect 368234 129574 368854 129658
rect 368234 129338 368266 129574
rect 368502 129338 368586 129574
rect 368822 129338 368854 129574
rect 368234 69894 368854 129338
rect 368234 69658 368266 69894
rect 368502 69658 368586 69894
rect 368822 69658 368854 69894
rect 368234 69574 368854 69658
rect 368234 69338 368266 69574
rect 368502 69338 368586 69574
rect 368822 69338 368854 69574
rect 368234 9894 368854 69338
rect 368234 9658 368266 9894
rect 368502 9658 368586 9894
rect 368822 9658 368854 9894
rect 368234 9574 368854 9658
rect 368234 9338 368266 9574
rect 368502 9338 368586 9574
rect 368822 9338 368854 9574
rect 368234 -4186 368854 9338
rect 368234 -4422 368266 -4186
rect 368502 -4422 368586 -4186
rect 368822 -4422 368854 -4186
rect 368234 -4506 368854 -4422
rect 368234 -4742 368266 -4506
rect 368502 -4742 368586 -4506
rect 368822 -4742 368854 -4506
rect 368234 -5734 368854 -4742
rect 371954 673614 372574 710042
rect 401954 711558 402574 711590
rect 401954 711322 401986 711558
rect 402222 711322 402306 711558
rect 402542 711322 402574 711558
rect 401954 711238 402574 711322
rect 401954 711002 401986 711238
rect 402222 711002 402306 711238
rect 402542 711002 402574 711238
rect 398234 709638 398854 709670
rect 398234 709402 398266 709638
rect 398502 709402 398586 709638
rect 398822 709402 398854 709638
rect 398234 709318 398854 709402
rect 398234 709082 398266 709318
rect 398502 709082 398586 709318
rect 398822 709082 398854 709318
rect 394514 707718 395134 707750
rect 394514 707482 394546 707718
rect 394782 707482 394866 707718
rect 395102 707482 395134 707718
rect 394514 707398 395134 707482
rect 394514 707162 394546 707398
rect 394782 707162 394866 707398
rect 395102 707162 395134 707398
rect 371954 673378 371986 673614
rect 372222 673378 372306 673614
rect 372542 673378 372574 673614
rect 371954 673294 372574 673378
rect 371954 673058 371986 673294
rect 372222 673058 372306 673294
rect 372542 673058 372574 673294
rect 371954 613614 372574 673058
rect 371954 613378 371986 613614
rect 372222 613378 372306 613614
rect 372542 613378 372574 613614
rect 371954 613294 372574 613378
rect 371954 613058 371986 613294
rect 372222 613058 372306 613294
rect 372542 613058 372574 613294
rect 371954 553614 372574 613058
rect 371954 553378 371986 553614
rect 372222 553378 372306 553614
rect 372542 553378 372574 553614
rect 371954 553294 372574 553378
rect 371954 553058 371986 553294
rect 372222 553058 372306 553294
rect 372542 553058 372574 553294
rect 371954 493614 372574 553058
rect 371954 493378 371986 493614
rect 372222 493378 372306 493614
rect 372542 493378 372574 493614
rect 371954 493294 372574 493378
rect 371954 493058 371986 493294
rect 372222 493058 372306 493294
rect 372542 493058 372574 493294
rect 371954 433614 372574 493058
rect 371954 433378 371986 433614
rect 372222 433378 372306 433614
rect 372542 433378 372574 433614
rect 371954 433294 372574 433378
rect 371954 433058 371986 433294
rect 372222 433058 372306 433294
rect 372542 433058 372574 433294
rect 371954 373614 372574 433058
rect 371954 373378 371986 373614
rect 372222 373378 372306 373614
rect 372542 373378 372574 373614
rect 371954 373294 372574 373378
rect 371954 373058 371986 373294
rect 372222 373058 372306 373294
rect 372542 373058 372574 373294
rect 371954 313614 372574 373058
rect 371954 313378 371986 313614
rect 372222 313378 372306 313614
rect 372542 313378 372574 313614
rect 371954 313294 372574 313378
rect 371954 313058 371986 313294
rect 372222 313058 372306 313294
rect 372542 313058 372574 313294
rect 371954 253614 372574 313058
rect 371954 253378 371986 253614
rect 372222 253378 372306 253614
rect 372542 253378 372574 253614
rect 371954 253294 372574 253378
rect 371954 253058 371986 253294
rect 372222 253058 372306 253294
rect 372542 253058 372574 253294
rect 371954 193614 372574 253058
rect 371954 193378 371986 193614
rect 372222 193378 372306 193614
rect 372542 193378 372574 193614
rect 371954 193294 372574 193378
rect 371954 193058 371986 193294
rect 372222 193058 372306 193294
rect 372542 193058 372574 193294
rect 371954 133614 372574 193058
rect 371954 133378 371986 133614
rect 372222 133378 372306 133614
rect 372542 133378 372574 133614
rect 371954 133294 372574 133378
rect 371954 133058 371986 133294
rect 372222 133058 372306 133294
rect 372542 133058 372574 133294
rect 371954 73614 372574 133058
rect 371954 73378 371986 73614
rect 372222 73378 372306 73614
rect 372542 73378 372574 73614
rect 371954 73294 372574 73378
rect 371954 73058 371986 73294
rect 372222 73058 372306 73294
rect 372542 73058 372574 73294
rect 371954 13614 372574 73058
rect 371954 13378 371986 13614
rect 372222 13378 372306 13614
rect 372542 13378 372574 13614
rect 371954 13294 372574 13378
rect 371954 13058 371986 13294
rect 372222 13058 372306 13294
rect 372542 13058 372574 13294
rect 341954 -7302 341986 -7066
rect 342222 -7302 342306 -7066
rect 342542 -7302 342574 -7066
rect 341954 -7386 342574 -7302
rect 341954 -7622 341986 -7386
rect 342222 -7622 342306 -7386
rect 342542 -7622 342574 -7386
rect 341954 -7654 342574 -7622
rect 371954 -6106 372574 13058
rect 390794 705798 391414 705830
rect 390794 705562 390826 705798
rect 391062 705562 391146 705798
rect 391382 705562 391414 705798
rect 390794 705478 391414 705562
rect 390794 705242 390826 705478
rect 391062 705242 391146 705478
rect 391382 705242 391414 705478
rect 390794 692454 391414 705242
rect 390794 692218 390826 692454
rect 391062 692218 391146 692454
rect 391382 692218 391414 692454
rect 390794 692134 391414 692218
rect 390794 691898 390826 692134
rect 391062 691898 391146 692134
rect 391382 691898 391414 692134
rect 390794 632454 391414 691898
rect 390794 632218 390826 632454
rect 391062 632218 391146 632454
rect 391382 632218 391414 632454
rect 390794 632134 391414 632218
rect 390794 631898 390826 632134
rect 391062 631898 391146 632134
rect 391382 631898 391414 632134
rect 390794 572454 391414 631898
rect 390794 572218 390826 572454
rect 391062 572218 391146 572454
rect 391382 572218 391414 572454
rect 390794 572134 391414 572218
rect 390794 571898 390826 572134
rect 391062 571898 391146 572134
rect 391382 571898 391414 572134
rect 390794 512454 391414 571898
rect 390794 512218 390826 512454
rect 391062 512218 391146 512454
rect 391382 512218 391414 512454
rect 390794 512134 391414 512218
rect 390794 511898 390826 512134
rect 391062 511898 391146 512134
rect 391382 511898 391414 512134
rect 390794 452454 391414 511898
rect 390794 452218 390826 452454
rect 391062 452218 391146 452454
rect 391382 452218 391414 452454
rect 390794 452134 391414 452218
rect 390794 451898 390826 452134
rect 391062 451898 391146 452134
rect 391382 451898 391414 452134
rect 390794 392454 391414 451898
rect 390794 392218 390826 392454
rect 391062 392218 391146 392454
rect 391382 392218 391414 392454
rect 390794 392134 391414 392218
rect 390794 391898 390826 392134
rect 391062 391898 391146 392134
rect 391382 391898 391414 392134
rect 390794 332454 391414 391898
rect 390794 332218 390826 332454
rect 391062 332218 391146 332454
rect 391382 332218 391414 332454
rect 390794 332134 391414 332218
rect 390794 331898 390826 332134
rect 391062 331898 391146 332134
rect 391382 331898 391414 332134
rect 390794 272454 391414 331898
rect 390794 272218 390826 272454
rect 391062 272218 391146 272454
rect 391382 272218 391414 272454
rect 390794 272134 391414 272218
rect 390794 271898 390826 272134
rect 391062 271898 391146 272134
rect 391382 271898 391414 272134
rect 390794 212454 391414 271898
rect 390794 212218 390826 212454
rect 391062 212218 391146 212454
rect 391382 212218 391414 212454
rect 390794 212134 391414 212218
rect 390794 211898 390826 212134
rect 391062 211898 391146 212134
rect 391382 211898 391414 212134
rect 390794 152454 391414 211898
rect 390794 152218 390826 152454
rect 391062 152218 391146 152454
rect 391382 152218 391414 152454
rect 390794 152134 391414 152218
rect 390794 151898 390826 152134
rect 391062 151898 391146 152134
rect 391382 151898 391414 152134
rect 390794 92454 391414 151898
rect 390794 92218 390826 92454
rect 391062 92218 391146 92454
rect 391382 92218 391414 92454
rect 390794 92134 391414 92218
rect 390794 91898 390826 92134
rect 391062 91898 391146 92134
rect 391382 91898 391414 92134
rect 390794 32454 391414 91898
rect 390794 32218 390826 32454
rect 391062 32218 391146 32454
rect 391382 32218 391414 32454
rect 390794 32134 391414 32218
rect 390794 31898 390826 32134
rect 391062 31898 391146 32134
rect 391382 31898 391414 32134
rect 390794 -1306 391414 31898
rect 390794 -1542 390826 -1306
rect 391062 -1542 391146 -1306
rect 391382 -1542 391414 -1306
rect 390794 -1626 391414 -1542
rect 390794 -1862 390826 -1626
rect 391062 -1862 391146 -1626
rect 391382 -1862 391414 -1626
rect 390794 -1894 391414 -1862
rect 394514 696174 395134 707162
rect 394514 695938 394546 696174
rect 394782 695938 394866 696174
rect 395102 695938 395134 696174
rect 394514 695854 395134 695938
rect 394514 695618 394546 695854
rect 394782 695618 394866 695854
rect 395102 695618 395134 695854
rect 394514 636174 395134 695618
rect 394514 635938 394546 636174
rect 394782 635938 394866 636174
rect 395102 635938 395134 636174
rect 394514 635854 395134 635938
rect 394514 635618 394546 635854
rect 394782 635618 394866 635854
rect 395102 635618 395134 635854
rect 394514 576174 395134 635618
rect 394514 575938 394546 576174
rect 394782 575938 394866 576174
rect 395102 575938 395134 576174
rect 394514 575854 395134 575938
rect 394514 575618 394546 575854
rect 394782 575618 394866 575854
rect 395102 575618 395134 575854
rect 394514 516174 395134 575618
rect 394514 515938 394546 516174
rect 394782 515938 394866 516174
rect 395102 515938 395134 516174
rect 394514 515854 395134 515938
rect 394514 515618 394546 515854
rect 394782 515618 394866 515854
rect 395102 515618 395134 515854
rect 394514 456174 395134 515618
rect 394514 455938 394546 456174
rect 394782 455938 394866 456174
rect 395102 455938 395134 456174
rect 394514 455854 395134 455938
rect 394514 455618 394546 455854
rect 394782 455618 394866 455854
rect 395102 455618 395134 455854
rect 394514 396174 395134 455618
rect 394514 395938 394546 396174
rect 394782 395938 394866 396174
rect 395102 395938 395134 396174
rect 394514 395854 395134 395938
rect 394514 395618 394546 395854
rect 394782 395618 394866 395854
rect 395102 395618 395134 395854
rect 394514 336174 395134 395618
rect 394514 335938 394546 336174
rect 394782 335938 394866 336174
rect 395102 335938 395134 336174
rect 394514 335854 395134 335938
rect 394514 335618 394546 335854
rect 394782 335618 394866 335854
rect 395102 335618 395134 335854
rect 394514 276174 395134 335618
rect 394514 275938 394546 276174
rect 394782 275938 394866 276174
rect 395102 275938 395134 276174
rect 394514 275854 395134 275938
rect 394514 275618 394546 275854
rect 394782 275618 394866 275854
rect 395102 275618 395134 275854
rect 394514 216174 395134 275618
rect 394514 215938 394546 216174
rect 394782 215938 394866 216174
rect 395102 215938 395134 216174
rect 394514 215854 395134 215938
rect 394514 215618 394546 215854
rect 394782 215618 394866 215854
rect 395102 215618 395134 215854
rect 394514 156174 395134 215618
rect 394514 155938 394546 156174
rect 394782 155938 394866 156174
rect 395102 155938 395134 156174
rect 394514 155854 395134 155938
rect 394514 155618 394546 155854
rect 394782 155618 394866 155854
rect 395102 155618 395134 155854
rect 394514 96174 395134 155618
rect 394514 95938 394546 96174
rect 394782 95938 394866 96174
rect 395102 95938 395134 96174
rect 394514 95854 395134 95938
rect 394514 95618 394546 95854
rect 394782 95618 394866 95854
rect 395102 95618 395134 95854
rect 394514 36174 395134 95618
rect 394514 35938 394546 36174
rect 394782 35938 394866 36174
rect 395102 35938 395134 36174
rect 394514 35854 395134 35938
rect 394514 35618 394546 35854
rect 394782 35618 394866 35854
rect 395102 35618 395134 35854
rect 394514 -3226 395134 35618
rect 394514 -3462 394546 -3226
rect 394782 -3462 394866 -3226
rect 395102 -3462 395134 -3226
rect 394514 -3546 395134 -3462
rect 394514 -3782 394546 -3546
rect 394782 -3782 394866 -3546
rect 395102 -3782 395134 -3546
rect 394514 -3814 395134 -3782
rect 398234 699894 398854 709082
rect 398234 699658 398266 699894
rect 398502 699658 398586 699894
rect 398822 699658 398854 699894
rect 398234 699574 398854 699658
rect 398234 699338 398266 699574
rect 398502 699338 398586 699574
rect 398822 699338 398854 699574
rect 398234 639894 398854 699338
rect 398234 639658 398266 639894
rect 398502 639658 398586 639894
rect 398822 639658 398854 639894
rect 398234 639574 398854 639658
rect 398234 639338 398266 639574
rect 398502 639338 398586 639574
rect 398822 639338 398854 639574
rect 398234 579894 398854 639338
rect 398234 579658 398266 579894
rect 398502 579658 398586 579894
rect 398822 579658 398854 579894
rect 398234 579574 398854 579658
rect 398234 579338 398266 579574
rect 398502 579338 398586 579574
rect 398822 579338 398854 579574
rect 398234 519894 398854 579338
rect 398234 519658 398266 519894
rect 398502 519658 398586 519894
rect 398822 519658 398854 519894
rect 398234 519574 398854 519658
rect 398234 519338 398266 519574
rect 398502 519338 398586 519574
rect 398822 519338 398854 519574
rect 398234 459894 398854 519338
rect 398234 459658 398266 459894
rect 398502 459658 398586 459894
rect 398822 459658 398854 459894
rect 398234 459574 398854 459658
rect 398234 459338 398266 459574
rect 398502 459338 398586 459574
rect 398822 459338 398854 459574
rect 398234 399894 398854 459338
rect 398234 399658 398266 399894
rect 398502 399658 398586 399894
rect 398822 399658 398854 399894
rect 398234 399574 398854 399658
rect 398234 399338 398266 399574
rect 398502 399338 398586 399574
rect 398822 399338 398854 399574
rect 398234 339894 398854 399338
rect 398234 339658 398266 339894
rect 398502 339658 398586 339894
rect 398822 339658 398854 339894
rect 398234 339574 398854 339658
rect 398234 339338 398266 339574
rect 398502 339338 398586 339574
rect 398822 339338 398854 339574
rect 398234 279894 398854 339338
rect 398234 279658 398266 279894
rect 398502 279658 398586 279894
rect 398822 279658 398854 279894
rect 398234 279574 398854 279658
rect 398234 279338 398266 279574
rect 398502 279338 398586 279574
rect 398822 279338 398854 279574
rect 398234 219894 398854 279338
rect 398234 219658 398266 219894
rect 398502 219658 398586 219894
rect 398822 219658 398854 219894
rect 398234 219574 398854 219658
rect 398234 219338 398266 219574
rect 398502 219338 398586 219574
rect 398822 219338 398854 219574
rect 398234 159894 398854 219338
rect 398234 159658 398266 159894
rect 398502 159658 398586 159894
rect 398822 159658 398854 159894
rect 398234 159574 398854 159658
rect 398234 159338 398266 159574
rect 398502 159338 398586 159574
rect 398822 159338 398854 159574
rect 398234 99894 398854 159338
rect 398234 99658 398266 99894
rect 398502 99658 398586 99894
rect 398822 99658 398854 99894
rect 398234 99574 398854 99658
rect 398234 99338 398266 99574
rect 398502 99338 398586 99574
rect 398822 99338 398854 99574
rect 398234 39894 398854 99338
rect 398234 39658 398266 39894
rect 398502 39658 398586 39894
rect 398822 39658 398854 39894
rect 398234 39574 398854 39658
rect 398234 39338 398266 39574
rect 398502 39338 398586 39574
rect 398822 39338 398854 39574
rect 398234 -5146 398854 39338
rect 398234 -5382 398266 -5146
rect 398502 -5382 398586 -5146
rect 398822 -5382 398854 -5146
rect 398234 -5466 398854 -5382
rect 398234 -5702 398266 -5466
rect 398502 -5702 398586 -5466
rect 398822 -5702 398854 -5466
rect 398234 -5734 398854 -5702
rect 401954 643614 402574 711002
rect 431954 710598 432574 711590
rect 431954 710362 431986 710598
rect 432222 710362 432306 710598
rect 432542 710362 432574 710598
rect 431954 710278 432574 710362
rect 431954 710042 431986 710278
rect 432222 710042 432306 710278
rect 432542 710042 432574 710278
rect 428234 708678 428854 709670
rect 428234 708442 428266 708678
rect 428502 708442 428586 708678
rect 428822 708442 428854 708678
rect 428234 708358 428854 708442
rect 428234 708122 428266 708358
rect 428502 708122 428586 708358
rect 428822 708122 428854 708358
rect 424514 706758 425134 707750
rect 424514 706522 424546 706758
rect 424782 706522 424866 706758
rect 425102 706522 425134 706758
rect 424514 706438 425134 706522
rect 424514 706202 424546 706438
rect 424782 706202 424866 706438
rect 425102 706202 425134 706438
rect 401954 643378 401986 643614
rect 402222 643378 402306 643614
rect 402542 643378 402574 643614
rect 401954 643294 402574 643378
rect 401954 643058 401986 643294
rect 402222 643058 402306 643294
rect 402542 643058 402574 643294
rect 401954 583614 402574 643058
rect 401954 583378 401986 583614
rect 402222 583378 402306 583614
rect 402542 583378 402574 583614
rect 401954 583294 402574 583378
rect 401954 583058 401986 583294
rect 402222 583058 402306 583294
rect 402542 583058 402574 583294
rect 401954 523614 402574 583058
rect 401954 523378 401986 523614
rect 402222 523378 402306 523614
rect 402542 523378 402574 523614
rect 401954 523294 402574 523378
rect 401954 523058 401986 523294
rect 402222 523058 402306 523294
rect 402542 523058 402574 523294
rect 401954 463614 402574 523058
rect 401954 463378 401986 463614
rect 402222 463378 402306 463614
rect 402542 463378 402574 463614
rect 401954 463294 402574 463378
rect 401954 463058 401986 463294
rect 402222 463058 402306 463294
rect 402542 463058 402574 463294
rect 401954 403614 402574 463058
rect 401954 403378 401986 403614
rect 402222 403378 402306 403614
rect 402542 403378 402574 403614
rect 401954 403294 402574 403378
rect 401954 403058 401986 403294
rect 402222 403058 402306 403294
rect 402542 403058 402574 403294
rect 401954 343614 402574 403058
rect 401954 343378 401986 343614
rect 402222 343378 402306 343614
rect 402542 343378 402574 343614
rect 401954 343294 402574 343378
rect 401954 343058 401986 343294
rect 402222 343058 402306 343294
rect 402542 343058 402574 343294
rect 401954 283614 402574 343058
rect 401954 283378 401986 283614
rect 402222 283378 402306 283614
rect 402542 283378 402574 283614
rect 401954 283294 402574 283378
rect 401954 283058 401986 283294
rect 402222 283058 402306 283294
rect 402542 283058 402574 283294
rect 401954 223614 402574 283058
rect 401954 223378 401986 223614
rect 402222 223378 402306 223614
rect 402542 223378 402574 223614
rect 401954 223294 402574 223378
rect 401954 223058 401986 223294
rect 402222 223058 402306 223294
rect 402542 223058 402574 223294
rect 401954 163614 402574 223058
rect 401954 163378 401986 163614
rect 402222 163378 402306 163614
rect 402542 163378 402574 163614
rect 401954 163294 402574 163378
rect 401954 163058 401986 163294
rect 402222 163058 402306 163294
rect 402542 163058 402574 163294
rect 401954 103614 402574 163058
rect 401954 103378 401986 103614
rect 402222 103378 402306 103614
rect 402542 103378 402574 103614
rect 401954 103294 402574 103378
rect 401954 103058 401986 103294
rect 402222 103058 402306 103294
rect 402542 103058 402574 103294
rect 401954 43614 402574 103058
rect 401954 43378 401986 43614
rect 402222 43378 402306 43614
rect 402542 43378 402574 43614
rect 401954 43294 402574 43378
rect 401954 43058 401986 43294
rect 402222 43058 402306 43294
rect 402542 43058 402574 43294
rect 371954 -6342 371986 -6106
rect 372222 -6342 372306 -6106
rect 372542 -6342 372574 -6106
rect 371954 -6426 372574 -6342
rect 371954 -6662 371986 -6426
rect 372222 -6662 372306 -6426
rect 372542 -6662 372574 -6426
rect 371954 -7654 372574 -6662
rect 401954 -7066 402574 43058
rect 420794 704838 421414 705830
rect 420794 704602 420826 704838
rect 421062 704602 421146 704838
rect 421382 704602 421414 704838
rect 420794 704518 421414 704602
rect 420794 704282 420826 704518
rect 421062 704282 421146 704518
rect 421382 704282 421414 704518
rect 420794 662454 421414 704282
rect 420794 662218 420826 662454
rect 421062 662218 421146 662454
rect 421382 662218 421414 662454
rect 420794 662134 421414 662218
rect 420794 661898 420826 662134
rect 421062 661898 421146 662134
rect 421382 661898 421414 662134
rect 420794 602454 421414 661898
rect 420794 602218 420826 602454
rect 421062 602218 421146 602454
rect 421382 602218 421414 602454
rect 420794 602134 421414 602218
rect 420794 601898 420826 602134
rect 421062 601898 421146 602134
rect 421382 601898 421414 602134
rect 420794 542454 421414 601898
rect 420794 542218 420826 542454
rect 421062 542218 421146 542454
rect 421382 542218 421414 542454
rect 420794 542134 421414 542218
rect 420794 541898 420826 542134
rect 421062 541898 421146 542134
rect 421382 541898 421414 542134
rect 420794 482454 421414 541898
rect 420794 482218 420826 482454
rect 421062 482218 421146 482454
rect 421382 482218 421414 482454
rect 420794 482134 421414 482218
rect 420794 481898 420826 482134
rect 421062 481898 421146 482134
rect 421382 481898 421414 482134
rect 420794 422454 421414 481898
rect 420794 422218 420826 422454
rect 421062 422218 421146 422454
rect 421382 422218 421414 422454
rect 420794 422134 421414 422218
rect 420794 421898 420826 422134
rect 421062 421898 421146 422134
rect 421382 421898 421414 422134
rect 420794 362454 421414 421898
rect 420794 362218 420826 362454
rect 421062 362218 421146 362454
rect 421382 362218 421414 362454
rect 420794 362134 421414 362218
rect 420794 361898 420826 362134
rect 421062 361898 421146 362134
rect 421382 361898 421414 362134
rect 420794 302454 421414 361898
rect 420794 302218 420826 302454
rect 421062 302218 421146 302454
rect 421382 302218 421414 302454
rect 420794 302134 421414 302218
rect 420794 301898 420826 302134
rect 421062 301898 421146 302134
rect 421382 301898 421414 302134
rect 420794 242454 421414 301898
rect 420794 242218 420826 242454
rect 421062 242218 421146 242454
rect 421382 242218 421414 242454
rect 420794 242134 421414 242218
rect 420794 241898 420826 242134
rect 421062 241898 421146 242134
rect 421382 241898 421414 242134
rect 420794 182454 421414 241898
rect 420794 182218 420826 182454
rect 421062 182218 421146 182454
rect 421382 182218 421414 182454
rect 420794 182134 421414 182218
rect 420794 181898 420826 182134
rect 421062 181898 421146 182134
rect 421382 181898 421414 182134
rect 420794 122454 421414 181898
rect 420794 122218 420826 122454
rect 421062 122218 421146 122454
rect 421382 122218 421414 122454
rect 420794 122134 421414 122218
rect 420794 121898 420826 122134
rect 421062 121898 421146 122134
rect 421382 121898 421414 122134
rect 420794 62454 421414 121898
rect 420794 62218 420826 62454
rect 421062 62218 421146 62454
rect 421382 62218 421414 62454
rect 420794 62134 421414 62218
rect 420794 61898 420826 62134
rect 421062 61898 421146 62134
rect 421382 61898 421414 62134
rect 420794 2454 421414 61898
rect 420794 2218 420826 2454
rect 421062 2218 421146 2454
rect 421382 2218 421414 2454
rect 420794 2134 421414 2218
rect 420794 1898 420826 2134
rect 421062 1898 421146 2134
rect 421382 1898 421414 2134
rect 420794 -346 421414 1898
rect 420794 -582 420826 -346
rect 421062 -582 421146 -346
rect 421382 -582 421414 -346
rect 420794 -666 421414 -582
rect 420794 -902 420826 -666
rect 421062 -902 421146 -666
rect 421382 -902 421414 -666
rect 420794 -1894 421414 -902
rect 424514 666174 425134 706202
rect 424514 665938 424546 666174
rect 424782 665938 424866 666174
rect 425102 665938 425134 666174
rect 424514 665854 425134 665938
rect 424514 665618 424546 665854
rect 424782 665618 424866 665854
rect 425102 665618 425134 665854
rect 424514 606174 425134 665618
rect 424514 605938 424546 606174
rect 424782 605938 424866 606174
rect 425102 605938 425134 606174
rect 424514 605854 425134 605938
rect 424514 605618 424546 605854
rect 424782 605618 424866 605854
rect 425102 605618 425134 605854
rect 424514 546174 425134 605618
rect 424514 545938 424546 546174
rect 424782 545938 424866 546174
rect 425102 545938 425134 546174
rect 424514 545854 425134 545938
rect 424514 545618 424546 545854
rect 424782 545618 424866 545854
rect 425102 545618 425134 545854
rect 424514 486174 425134 545618
rect 424514 485938 424546 486174
rect 424782 485938 424866 486174
rect 425102 485938 425134 486174
rect 424514 485854 425134 485938
rect 424514 485618 424546 485854
rect 424782 485618 424866 485854
rect 425102 485618 425134 485854
rect 424514 426174 425134 485618
rect 424514 425938 424546 426174
rect 424782 425938 424866 426174
rect 425102 425938 425134 426174
rect 424514 425854 425134 425938
rect 424514 425618 424546 425854
rect 424782 425618 424866 425854
rect 425102 425618 425134 425854
rect 424514 366174 425134 425618
rect 424514 365938 424546 366174
rect 424782 365938 424866 366174
rect 425102 365938 425134 366174
rect 424514 365854 425134 365938
rect 424514 365618 424546 365854
rect 424782 365618 424866 365854
rect 425102 365618 425134 365854
rect 424514 306174 425134 365618
rect 424514 305938 424546 306174
rect 424782 305938 424866 306174
rect 425102 305938 425134 306174
rect 424514 305854 425134 305938
rect 424514 305618 424546 305854
rect 424782 305618 424866 305854
rect 425102 305618 425134 305854
rect 424514 246174 425134 305618
rect 424514 245938 424546 246174
rect 424782 245938 424866 246174
rect 425102 245938 425134 246174
rect 424514 245854 425134 245938
rect 424514 245618 424546 245854
rect 424782 245618 424866 245854
rect 425102 245618 425134 245854
rect 424514 186174 425134 245618
rect 424514 185938 424546 186174
rect 424782 185938 424866 186174
rect 425102 185938 425134 186174
rect 424514 185854 425134 185938
rect 424514 185618 424546 185854
rect 424782 185618 424866 185854
rect 425102 185618 425134 185854
rect 424514 126174 425134 185618
rect 424514 125938 424546 126174
rect 424782 125938 424866 126174
rect 425102 125938 425134 126174
rect 424514 125854 425134 125938
rect 424514 125618 424546 125854
rect 424782 125618 424866 125854
rect 425102 125618 425134 125854
rect 424514 66174 425134 125618
rect 424514 65938 424546 66174
rect 424782 65938 424866 66174
rect 425102 65938 425134 66174
rect 424514 65854 425134 65938
rect 424514 65618 424546 65854
rect 424782 65618 424866 65854
rect 425102 65618 425134 65854
rect 424514 6174 425134 65618
rect 424514 5938 424546 6174
rect 424782 5938 424866 6174
rect 425102 5938 425134 6174
rect 424514 5854 425134 5938
rect 424514 5618 424546 5854
rect 424782 5618 424866 5854
rect 425102 5618 425134 5854
rect 424514 -2266 425134 5618
rect 424514 -2502 424546 -2266
rect 424782 -2502 424866 -2266
rect 425102 -2502 425134 -2266
rect 424514 -2586 425134 -2502
rect 424514 -2822 424546 -2586
rect 424782 -2822 424866 -2586
rect 425102 -2822 425134 -2586
rect 424514 -3814 425134 -2822
rect 428234 669894 428854 708122
rect 428234 669658 428266 669894
rect 428502 669658 428586 669894
rect 428822 669658 428854 669894
rect 428234 669574 428854 669658
rect 428234 669338 428266 669574
rect 428502 669338 428586 669574
rect 428822 669338 428854 669574
rect 428234 609894 428854 669338
rect 428234 609658 428266 609894
rect 428502 609658 428586 609894
rect 428822 609658 428854 609894
rect 428234 609574 428854 609658
rect 428234 609338 428266 609574
rect 428502 609338 428586 609574
rect 428822 609338 428854 609574
rect 428234 549894 428854 609338
rect 428234 549658 428266 549894
rect 428502 549658 428586 549894
rect 428822 549658 428854 549894
rect 428234 549574 428854 549658
rect 428234 549338 428266 549574
rect 428502 549338 428586 549574
rect 428822 549338 428854 549574
rect 428234 489894 428854 549338
rect 428234 489658 428266 489894
rect 428502 489658 428586 489894
rect 428822 489658 428854 489894
rect 428234 489574 428854 489658
rect 428234 489338 428266 489574
rect 428502 489338 428586 489574
rect 428822 489338 428854 489574
rect 428234 429894 428854 489338
rect 428234 429658 428266 429894
rect 428502 429658 428586 429894
rect 428822 429658 428854 429894
rect 428234 429574 428854 429658
rect 428234 429338 428266 429574
rect 428502 429338 428586 429574
rect 428822 429338 428854 429574
rect 428234 369894 428854 429338
rect 428234 369658 428266 369894
rect 428502 369658 428586 369894
rect 428822 369658 428854 369894
rect 428234 369574 428854 369658
rect 428234 369338 428266 369574
rect 428502 369338 428586 369574
rect 428822 369338 428854 369574
rect 428234 309894 428854 369338
rect 428234 309658 428266 309894
rect 428502 309658 428586 309894
rect 428822 309658 428854 309894
rect 428234 309574 428854 309658
rect 428234 309338 428266 309574
rect 428502 309338 428586 309574
rect 428822 309338 428854 309574
rect 428234 249894 428854 309338
rect 428234 249658 428266 249894
rect 428502 249658 428586 249894
rect 428822 249658 428854 249894
rect 428234 249574 428854 249658
rect 428234 249338 428266 249574
rect 428502 249338 428586 249574
rect 428822 249338 428854 249574
rect 428234 189894 428854 249338
rect 428234 189658 428266 189894
rect 428502 189658 428586 189894
rect 428822 189658 428854 189894
rect 428234 189574 428854 189658
rect 428234 189338 428266 189574
rect 428502 189338 428586 189574
rect 428822 189338 428854 189574
rect 428234 129894 428854 189338
rect 428234 129658 428266 129894
rect 428502 129658 428586 129894
rect 428822 129658 428854 129894
rect 428234 129574 428854 129658
rect 428234 129338 428266 129574
rect 428502 129338 428586 129574
rect 428822 129338 428854 129574
rect 428234 69894 428854 129338
rect 428234 69658 428266 69894
rect 428502 69658 428586 69894
rect 428822 69658 428854 69894
rect 428234 69574 428854 69658
rect 428234 69338 428266 69574
rect 428502 69338 428586 69574
rect 428822 69338 428854 69574
rect 428234 9894 428854 69338
rect 428234 9658 428266 9894
rect 428502 9658 428586 9894
rect 428822 9658 428854 9894
rect 428234 9574 428854 9658
rect 428234 9338 428266 9574
rect 428502 9338 428586 9574
rect 428822 9338 428854 9574
rect 428234 -4186 428854 9338
rect 428234 -4422 428266 -4186
rect 428502 -4422 428586 -4186
rect 428822 -4422 428854 -4186
rect 428234 -4506 428854 -4422
rect 428234 -4742 428266 -4506
rect 428502 -4742 428586 -4506
rect 428822 -4742 428854 -4506
rect 428234 -5734 428854 -4742
rect 431954 673614 432574 710042
rect 461954 711558 462574 711590
rect 461954 711322 461986 711558
rect 462222 711322 462306 711558
rect 462542 711322 462574 711558
rect 461954 711238 462574 711322
rect 461954 711002 461986 711238
rect 462222 711002 462306 711238
rect 462542 711002 462574 711238
rect 458234 709638 458854 709670
rect 458234 709402 458266 709638
rect 458502 709402 458586 709638
rect 458822 709402 458854 709638
rect 458234 709318 458854 709402
rect 458234 709082 458266 709318
rect 458502 709082 458586 709318
rect 458822 709082 458854 709318
rect 454514 707718 455134 707750
rect 454514 707482 454546 707718
rect 454782 707482 454866 707718
rect 455102 707482 455134 707718
rect 454514 707398 455134 707482
rect 454514 707162 454546 707398
rect 454782 707162 454866 707398
rect 455102 707162 455134 707398
rect 431954 673378 431986 673614
rect 432222 673378 432306 673614
rect 432542 673378 432574 673614
rect 431954 673294 432574 673378
rect 431954 673058 431986 673294
rect 432222 673058 432306 673294
rect 432542 673058 432574 673294
rect 431954 613614 432574 673058
rect 431954 613378 431986 613614
rect 432222 613378 432306 613614
rect 432542 613378 432574 613614
rect 431954 613294 432574 613378
rect 431954 613058 431986 613294
rect 432222 613058 432306 613294
rect 432542 613058 432574 613294
rect 431954 553614 432574 613058
rect 431954 553378 431986 553614
rect 432222 553378 432306 553614
rect 432542 553378 432574 553614
rect 431954 553294 432574 553378
rect 431954 553058 431986 553294
rect 432222 553058 432306 553294
rect 432542 553058 432574 553294
rect 431954 493614 432574 553058
rect 431954 493378 431986 493614
rect 432222 493378 432306 493614
rect 432542 493378 432574 493614
rect 431954 493294 432574 493378
rect 431954 493058 431986 493294
rect 432222 493058 432306 493294
rect 432542 493058 432574 493294
rect 431954 433614 432574 493058
rect 431954 433378 431986 433614
rect 432222 433378 432306 433614
rect 432542 433378 432574 433614
rect 431954 433294 432574 433378
rect 431954 433058 431986 433294
rect 432222 433058 432306 433294
rect 432542 433058 432574 433294
rect 431954 373614 432574 433058
rect 431954 373378 431986 373614
rect 432222 373378 432306 373614
rect 432542 373378 432574 373614
rect 431954 373294 432574 373378
rect 431954 373058 431986 373294
rect 432222 373058 432306 373294
rect 432542 373058 432574 373294
rect 431954 313614 432574 373058
rect 431954 313378 431986 313614
rect 432222 313378 432306 313614
rect 432542 313378 432574 313614
rect 431954 313294 432574 313378
rect 431954 313058 431986 313294
rect 432222 313058 432306 313294
rect 432542 313058 432574 313294
rect 431954 253614 432574 313058
rect 431954 253378 431986 253614
rect 432222 253378 432306 253614
rect 432542 253378 432574 253614
rect 431954 253294 432574 253378
rect 431954 253058 431986 253294
rect 432222 253058 432306 253294
rect 432542 253058 432574 253294
rect 431954 193614 432574 253058
rect 431954 193378 431986 193614
rect 432222 193378 432306 193614
rect 432542 193378 432574 193614
rect 431954 193294 432574 193378
rect 431954 193058 431986 193294
rect 432222 193058 432306 193294
rect 432542 193058 432574 193294
rect 431954 133614 432574 193058
rect 431954 133378 431986 133614
rect 432222 133378 432306 133614
rect 432542 133378 432574 133614
rect 431954 133294 432574 133378
rect 431954 133058 431986 133294
rect 432222 133058 432306 133294
rect 432542 133058 432574 133294
rect 431954 73614 432574 133058
rect 431954 73378 431986 73614
rect 432222 73378 432306 73614
rect 432542 73378 432574 73614
rect 431954 73294 432574 73378
rect 431954 73058 431986 73294
rect 432222 73058 432306 73294
rect 432542 73058 432574 73294
rect 431954 13614 432574 73058
rect 431954 13378 431986 13614
rect 432222 13378 432306 13614
rect 432542 13378 432574 13614
rect 431954 13294 432574 13378
rect 431954 13058 431986 13294
rect 432222 13058 432306 13294
rect 432542 13058 432574 13294
rect 401954 -7302 401986 -7066
rect 402222 -7302 402306 -7066
rect 402542 -7302 402574 -7066
rect 401954 -7386 402574 -7302
rect 401954 -7622 401986 -7386
rect 402222 -7622 402306 -7386
rect 402542 -7622 402574 -7386
rect 401954 -7654 402574 -7622
rect 431954 -6106 432574 13058
rect 450794 705798 451414 705830
rect 450794 705562 450826 705798
rect 451062 705562 451146 705798
rect 451382 705562 451414 705798
rect 450794 705478 451414 705562
rect 450794 705242 450826 705478
rect 451062 705242 451146 705478
rect 451382 705242 451414 705478
rect 450794 692454 451414 705242
rect 450794 692218 450826 692454
rect 451062 692218 451146 692454
rect 451382 692218 451414 692454
rect 450794 692134 451414 692218
rect 450794 691898 450826 692134
rect 451062 691898 451146 692134
rect 451382 691898 451414 692134
rect 450794 632454 451414 691898
rect 450794 632218 450826 632454
rect 451062 632218 451146 632454
rect 451382 632218 451414 632454
rect 450794 632134 451414 632218
rect 450794 631898 450826 632134
rect 451062 631898 451146 632134
rect 451382 631898 451414 632134
rect 450794 572454 451414 631898
rect 450794 572218 450826 572454
rect 451062 572218 451146 572454
rect 451382 572218 451414 572454
rect 450794 572134 451414 572218
rect 450794 571898 450826 572134
rect 451062 571898 451146 572134
rect 451382 571898 451414 572134
rect 450794 512454 451414 571898
rect 450794 512218 450826 512454
rect 451062 512218 451146 512454
rect 451382 512218 451414 512454
rect 450794 512134 451414 512218
rect 450794 511898 450826 512134
rect 451062 511898 451146 512134
rect 451382 511898 451414 512134
rect 450794 452454 451414 511898
rect 450794 452218 450826 452454
rect 451062 452218 451146 452454
rect 451382 452218 451414 452454
rect 450794 452134 451414 452218
rect 450794 451898 450826 452134
rect 451062 451898 451146 452134
rect 451382 451898 451414 452134
rect 450794 392454 451414 451898
rect 450794 392218 450826 392454
rect 451062 392218 451146 392454
rect 451382 392218 451414 392454
rect 450794 392134 451414 392218
rect 450794 391898 450826 392134
rect 451062 391898 451146 392134
rect 451382 391898 451414 392134
rect 450794 332454 451414 391898
rect 450794 332218 450826 332454
rect 451062 332218 451146 332454
rect 451382 332218 451414 332454
rect 450794 332134 451414 332218
rect 450794 331898 450826 332134
rect 451062 331898 451146 332134
rect 451382 331898 451414 332134
rect 450794 272454 451414 331898
rect 450794 272218 450826 272454
rect 451062 272218 451146 272454
rect 451382 272218 451414 272454
rect 450794 272134 451414 272218
rect 450794 271898 450826 272134
rect 451062 271898 451146 272134
rect 451382 271898 451414 272134
rect 450794 212454 451414 271898
rect 450794 212218 450826 212454
rect 451062 212218 451146 212454
rect 451382 212218 451414 212454
rect 450794 212134 451414 212218
rect 450794 211898 450826 212134
rect 451062 211898 451146 212134
rect 451382 211898 451414 212134
rect 450794 152454 451414 211898
rect 450794 152218 450826 152454
rect 451062 152218 451146 152454
rect 451382 152218 451414 152454
rect 450794 152134 451414 152218
rect 450794 151898 450826 152134
rect 451062 151898 451146 152134
rect 451382 151898 451414 152134
rect 450794 92454 451414 151898
rect 450794 92218 450826 92454
rect 451062 92218 451146 92454
rect 451382 92218 451414 92454
rect 450794 92134 451414 92218
rect 450794 91898 450826 92134
rect 451062 91898 451146 92134
rect 451382 91898 451414 92134
rect 450794 32454 451414 91898
rect 450794 32218 450826 32454
rect 451062 32218 451146 32454
rect 451382 32218 451414 32454
rect 450794 32134 451414 32218
rect 450794 31898 450826 32134
rect 451062 31898 451146 32134
rect 451382 31898 451414 32134
rect 450794 -1306 451414 31898
rect 450794 -1542 450826 -1306
rect 451062 -1542 451146 -1306
rect 451382 -1542 451414 -1306
rect 450794 -1626 451414 -1542
rect 450794 -1862 450826 -1626
rect 451062 -1862 451146 -1626
rect 451382 -1862 451414 -1626
rect 450794 -1894 451414 -1862
rect 454514 696174 455134 707162
rect 454514 695938 454546 696174
rect 454782 695938 454866 696174
rect 455102 695938 455134 696174
rect 454514 695854 455134 695938
rect 454514 695618 454546 695854
rect 454782 695618 454866 695854
rect 455102 695618 455134 695854
rect 454514 636174 455134 695618
rect 454514 635938 454546 636174
rect 454782 635938 454866 636174
rect 455102 635938 455134 636174
rect 454514 635854 455134 635938
rect 454514 635618 454546 635854
rect 454782 635618 454866 635854
rect 455102 635618 455134 635854
rect 454514 576174 455134 635618
rect 454514 575938 454546 576174
rect 454782 575938 454866 576174
rect 455102 575938 455134 576174
rect 454514 575854 455134 575938
rect 454514 575618 454546 575854
rect 454782 575618 454866 575854
rect 455102 575618 455134 575854
rect 454514 516174 455134 575618
rect 454514 515938 454546 516174
rect 454782 515938 454866 516174
rect 455102 515938 455134 516174
rect 454514 515854 455134 515938
rect 454514 515618 454546 515854
rect 454782 515618 454866 515854
rect 455102 515618 455134 515854
rect 454514 456174 455134 515618
rect 454514 455938 454546 456174
rect 454782 455938 454866 456174
rect 455102 455938 455134 456174
rect 454514 455854 455134 455938
rect 454514 455618 454546 455854
rect 454782 455618 454866 455854
rect 455102 455618 455134 455854
rect 454514 396174 455134 455618
rect 454514 395938 454546 396174
rect 454782 395938 454866 396174
rect 455102 395938 455134 396174
rect 454514 395854 455134 395938
rect 454514 395618 454546 395854
rect 454782 395618 454866 395854
rect 455102 395618 455134 395854
rect 454514 336174 455134 395618
rect 454514 335938 454546 336174
rect 454782 335938 454866 336174
rect 455102 335938 455134 336174
rect 454514 335854 455134 335938
rect 454514 335618 454546 335854
rect 454782 335618 454866 335854
rect 455102 335618 455134 335854
rect 454514 276174 455134 335618
rect 454514 275938 454546 276174
rect 454782 275938 454866 276174
rect 455102 275938 455134 276174
rect 454514 275854 455134 275938
rect 454514 275618 454546 275854
rect 454782 275618 454866 275854
rect 455102 275618 455134 275854
rect 454514 216174 455134 275618
rect 454514 215938 454546 216174
rect 454782 215938 454866 216174
rect 455102 215938 455134 216174
rect 454514 215854 455134 215938
rect 454514 215618 454546 215854
rect 454782 215618 454866 215854
rect 455102 215618 455134 215854
rect 454514 156174 455134 215618
rect 454514 155938 454546 156174
rect 454782 155938 454866 156174
rect 455102 155938 455134 156174
rect 454514 155854 455134 155938
rect 454514 155618 454546 155854
rect 454782 155618 454866 155854
rect 455102 155618 455134 155854
rect 454514 96174 455134 155618
rect 454514 95938 454546 96174
rect 454782 95938 454866 96174
rect 455102 95938 455134 96174
rect 454514 95854 455134 95938
rect 454514 95618 454546 95854
rect 454782 95618 454866 95854
rect 455102 95618 455134 95854
rect 454514 36174 455134 95618
rect 454514 35938 454546 36174
rect 454782 35938 454866 36174
rect 455102 35938 455134 36174
rect 454514 35854 455134 35938
rect 454514 35618 454546 35854
rect 454782 35618 454866 35854
rect 455102 35618 455134 35854
rect 454514 -3226 455134 35618
rect 454514 -3462 454546 -3226
rect 454782 -3462 454866 -3226
rect 455102 -3462 455134 -3226
rect 454514 -3546 455134 -3462
rect 454514 -3782 454546 -3546
rect 454782 -3782 454866 -3546
rect 455102 -3782 455134 -3546
rect 454514 -3814 455134 -3782
rect 458234 699894 458854 709082
rect 458234 699658 458266 699894
rect 458502 699658 458586 699894
rect 458822 699658 458854 699894
rect 458234 699574 458854 699658
rect 458234 699338 458266 699574
rect 458502 699338 458586 699574
rect 458822 699338 458854 699574
rect 458234 639894 458854 699338
rect 458234 639658 458266 639894
rect 458502 639658 458586 639894
rect 458822 639658 458854 639894
rect 458234 639574 458854 639658
rect 458234 639338 458266 639574
rect 458502 639338 458586 639574
rect 458822 639338 458854 639574
rect 458234 579894 458854 639338
rect 458234 579658 458266 579894
rect 458502 579658 458586 579894
rect 458822 579658 458854 579894
rect 458234 579574 458854 579658
rect 458234 579338 458266 579574
rect 458502 579338 458586 579574
rect 458822 579338 458854 579574
rect 458234 519894 458854 579338
rect 458234 519658 458266 519894
rect 458502 519658 458586 519894
rect 458822 519658 458854 519894
rect 458234 519574 458854 519658
rect 458234 519338 458266 519574
rect 458502 519338 458586 519574
rect 458822 519338 458854 519574
rect 458234 459894 458854 519338
rect 458234 459658 458266 459894
rect 458502 459658 458586 459894
rect 458822 459658 458854 459894
rect 458234 459574 458854 459658
rect 458234 459338 458266 459574
rect 458502 459338 458586 459574
rect 458822 459338 458854 459574
rect 458234 399894 458854 459338
rect 458234 399658 458266 399894
rect 458502 399658 458586 399894
rect 458822 399658 458854 399894
rect 458234 399574 458854 399658
rect 458234 399338 458266 399574
rect 458502 399338 458586 399574
rect 458822 399338 458854 399574
rect 458234 339894 458854 399338
rect 458234 339658 458266 339894
rect 458502 339658 458586 339894
rect 458822 339658 458854 339894
rect 458234 339574 458854 339658
rect 458234 339338 458266 339574
rect 458502 339338 458586 339574
rect 458822 339338 458854 339574
rect 458234 279894 458854 339338
rect 458234 279658 458266 279894
rect 458502 279658 458586 279894
rect 458822 279658 458854 279894
rect 458234 279574 458854 279658
rect 458234 279338 458266 279574
rect 458502 279338 458586 279574
rect 458822 279338 458854 279574
rect 458234 219894 458854 279338
rect 458234 219658 458266 219894
rect 458502 219658 458586 219894
rect 458822 219658 458854 219894
rect 458234 219574 458854 219658
rect 458234 219338 458266 219574
rect 458502 219338 458586 219574
rect 458822 219338 458854 219574
rect 458234 159894 458854 219338
rect 458234 159658 458266 159894
rect 458502 159658 458586 159894
rect 458822 159658 458854 159894
rect 458234 159574 458854 159658
rect 458234 159338 458266 159574
rect 458502 159338 458586 159574
rect 458822 159338 458854 159574
rect 458234 99894 458854 159338
rect 458234 99658 458266 99894
rect 458502 99658 458586 99894
rect 458822 99658 458854 99894
rect 458234 99574 458854 99658
rect 458234 99338 458266 99574
rect 458502 99338 458586 99574
rect 458822 99338 458854 99574
rect 458234 39894 458854 99338
rect 458234 39658 458266 39894
rect 458502 39658 458586 39894
rect 458822 39658 458854 39894
rect 458234 39574 458854 39658
rect 458234 39338 458266 39574
rect 458502 39338 458586 39574
rect 458822 39338 458854 39574
rect 458234 -5146 458854 39338
rect 458234 -5382 458266 -5146
rect 458502 -5382 458586 -5146
rect 458822 -5382 458854 -5146
rect 458234 -5466 458854 -5382
rect 458234 -5702 458266 -5466
rect 458502 -5702 458586 -5466
rect 458822 -5702 458854 -5466
rect 458234 -5734 458854 -5702
rect 461954 643614 462574 711002
rect 491954 710598 492574 711590
rect 491954 710362 491986 710598
rect 492222 710362 492306 710598
rect 492542 710362 492574 710598
rect 491954 710278 492574 710362
rect 491954 710042 491986 710278
rect 492222 710042 492306 710278
rect 492542 710042 492574 710278
rect 488234 708678 488854 709670
rect 488234 708442 488266 708678
rect 488502 708442 488586 708678
rect 488822 708442 488854 708678
rect 488234 708358 488854 708442
rect 488234 708122 488266 708358
rect 488502 708122 488586 708358
rect 488822 708122 488854 708358
rect 484514 706758 485134 707750
rect 484514 706522 484546 706758
rect 484782 706522 484866 706758
rect 485102 706522 485134 706758
rect 484514 706438 485134 706522
rect 484514 706202 484546 706438
rect 484782 706202 484866 706438
rect 485102 706202 485134 706438
rect 461954 643378 461986 643614
rect 462222 643378 462306 643614
rect 462542 643378 462574 643614
rect 461954 643294 462574 643378
rect 461954 643058 461986 643294
rect 462222 643058 462306 643294
rect 462542 643058 462574 643294
rect 461954 583614 462574 643058
rect 461954 583378 461986 583614
rect 462222 583378 462306 583614
rect 462542 583378 462574 583614
rect 461954 583294 462574 583378
rect 461954 583058 461986 583294
rect 462222 583058 462306 583294
rect 462542 583058 462574 583294
rect 461954 523614 462574 583058
rect 461954 523378 461986 523614
rect 462222 523378 462306 523614
rect 462542 523378 462574 523614
rect 461954 523294 462574 523378
rect 461954 523058 461986 523294
rect 462222 523058 462306 523294
rect 462542 523058 462574 523294
rect 461954 463614 462574 523058
rect 461954 463378 461986 463614
rect 462222 463378 462306 463614
rect 462542 463378 462574 463614
rect 461954 463294 462574 463378
rect 461954 463058 461986 463294
rect 462222 463058 462306 463294
rect 462542 463058 462574 463294
rect 461954 403614 462574 463058
rect 461954 403378 461986 403614
rect 462222 403378 462306 403614
rect 462542 403378 462574 403614
rect 461954 403294 462574 403378
rect 461954 403058 461986 403294
rect 462222 403058 462306 403294
rect 462542 403058 462574 403294
rect 461954 343614 462574 403058
rect 461954 343378 461986 343614
rect 462222 343378 462306 343614
rect 462542 343378 462574 343614
rect 461954 343294 462574 343378
rect 461954 343058 461986 343294
rect 462222 343058 462306 343294
rect 462542 343058 462574 343294
rect 461954 283614 462574 343058
rect 461954 283378 461986 283614
rect 462222 283378 462306 283614
rect 462542 283378 462574 283614
rect 461954 283294 462574 283378
rect 461954 283058 461986 283294
rect 462222 283058 462306 283294
rect 462542 283058 462574 283294
rect 461954 223614 462574 283058
rect 461954 223378 461986 223614
rect 462222 223378 462306 223614
rect 462542 223378 462574 223614
rect 461954 223294 462574 223378
rect 461954 223058 461986 223294
rect 462222 223058 462306 223294
rect 462542 223058 462574 223294
rect 461954 163614 462574 223058
rect 461954 163378 461986 163614
rect 462222 163378 462306 163614
rect 462542 163378 462574 163614
rect 461954 163294 462574 163378
rect 461954 163058 461986 163294
rect 462222 163058 462306 163294
rect 462542 163058 462574 163294
rect 461954 103614 462574 163058
rect 461954 103378 461986 103614
rect 462222 103378 462306 103614
rect 462542 103378 462574 103614
rect 461954 103294 462574 103378
rect 461954 103058 461986 103294
rect 462222 103058 462306 103294
rect 462542 103058 462574 103294
rect 461954 43614 462574 103058
rect 461954 43378 461986 43614
rect 462222 43378 462306 43614
rect 462542 43378 462574 43614
rect 461954 43294 462574 43378
rect 461954 43058 461986 43294
rect 462222 43058 462306 43294
rect 462542 43058 462574 43294
rect 431954 -6342 431986 -6106
rect 432222 -6342 432306 -6106
rect 432542 -6342 432574 -6106
rect 431954 -6426 432574 -6342
rect 431954 -6662 431986 -6426
rect 432222 -6662 432306 -6426
rect 432542 -6662 432574 -6426
rect 431954 -7654 432574 -6662
rect 461954 -7066 462574 43058
rect 480794 704838 481414 705830
rect 480794 704602 480826 704838
rect 481062 704602 481146 704838
rect 481382 704602 481414 704838
rect 480794 704518 481414 704602
rect 480794 704282 480826 704518
rect 481062 704282 481146 704518
rect 481382 704282 481414 704518
rect 480794 662454 481414 704282
rect 480794 662218 480826 662454
rect 481062 662218 481146 662454
rect 481382 662218 481414 662454
rect 480794 662134 481414 662218
rect 480794 661898 480826 662134
rect 481062 661898 481146 662134
rect 481382 661898 481414 662134
rect 480794 602454 481414 661898
rect 480794 602218 480826 602454
rect 481062 602218 481146 602454
rect 481382 602218 481414 602454
rect 480794 602134 481414 602218
rect 480794 601898 480826 602134
rect 481062 601898 481146 602134
rect 481382 601898 481414 602134
rect 480794 542454 481414 601898
rect 480794 542218 480826 542454
rect 481062 542218 481146 542454
rect 481382 542218 481414 542454
rect 480794 542134 481414 542218
rect 480794 541898 480826 542134
rect 481062 541898 481146 542134
rect 481382 541898 481414 542134
rect 480794 482454 481414 541898
rect 480794 482218 480826 482454
rect 481062 482218 481146 482454
rect 481382 482218 481414 482454
rect 480794 482134 481414 482218
rect 480794 481898 480826 482134
rect 481062 481898 481146 482134
rect 481382 481898 481414 482134
rect 480794 422454 481414 481898
rect 480794 422218 480826 422454
rect 481062 422218 481146 422454
rect 481382 422218 481414 422454
rect 480794 422134 481414 422218
rect 480794 421898 480826 422134
rect 481062 421898 481146 422134
rect 481382 421898 481414 422134
rect 480794 362454 481414 421898
rect 480794 362218 480826 362454
rect 481062 362218 481146 362454
rect 481382 362218 481414 362454
rect 480794 362134 481414 362218
rect 480794 361898 480826 362134
rect 481062 361898 481146 362134
rect 481382 361898 481414 362134
rect 480794 302454 481414 361898
rect 480794 302218 480826 302454
rect 481062 302218 481146 302454
rect 481382 302218 481414 302454
rect 480794 302134 481414 302218
rect 480794 301898 480826 302134
rect 481062 301898 481146 302134
rect 481382 301898 481414 302134
rect 480794 242454 481414 301898
rect 480794 242218 480826 242454
rect 481062 242218 481146 242454
rect 481382 242218 481414 242454
rect 480794 242134 481414 242218
rect 480794 241898 480826 242134
rect 481062 241898 481146 242134
rect 481382 241898 481414 242134
rect 480794 182454 481414 241898
rect 480794 182218 480826 182454
rect 481062 182218 481146 182454
rect 481382 182218 481414 182454
rect 480794 182134 481414 182218
rect 480794 181898 480826 182134
rect 481062 181898 481146 182134
rect 481382 181898 481414 182134
rect 480794 122454 481414 181898
rect 480794 122218 480826 122454
rect 481062 122218 481146 122454
rect 481382 122218 481414 122454
rect 480794 122134 481414 122218
rect 480794 121898 480826 122134
rect 481062 121898 481146 122134
rect 481382 121898 481414 122134
rect 480794 62454 481414 121898
rect 480794 62218 480826 62454
rect 481062 62218 481146 62454
rect 481382 62218 481414 62454
rect 480794 62134 481414 62218
rect 480794 61898 480826 62134
rect 481062 61898 481146 62134
rect 481382 61898 481414 62134
rect 480794 2454 481414 61898
rect 480794 2218 480826 2454
rect 481062 2218 481146 2454
rect 481382 2218 481414 2454
rect 480794 2134 481414 2218
rect 480794 1898 480826 2134
rect 481062 1898 481146 2134
rect 481382 1898 481414 2134
rect 480794 -346 481414 1898
rect 480794 -582 480826 -346
rect 481062 -582 481146 -346
rect 481382 -582 481414 -346
rect 480794 -666 481414 -582
rect 480794 -902 480826 -666
rect 481062 -902 481146 -666
rect 481382 -902 481414 -666
rect 480794 -1894 481414 -902
rect 484514 666174 485134 706202
rect 484514 665938 484546 666174
rect 484782 665938 484866 666174
rect 485102 665938 485134 666174
rect 484514 665854 485134 665938
rect 484514 665618 484546 665854
rect 484782 665618 484866 665854
rect 485102 665618 485134 665854
rect 484514 606174 485134 665618
rect 484514 605938 484546 606174
rect 484782 605938 484866 606174
rect 485102 605938 485134 606174
rect 484514 605854 485134 605938
rect 484514 605618 484546 605854
rect 484782 605618 484866 605854
rect 485102 605618 485134 605854
rect 484514 546174 485134 605618
rect 484514 545938 484546 546174
rect 484782 545938 484866 546174
rect 485102 545938 485134 546174
rect 484514 545854 485134 545938
rect 484514 545618 484546 545854
rect 484782 545618 484866 545854
rect 485102 545618 485134 545854
rect 484514 486174 485134 545618
rect 484514 485938 484546 486174
rect 484782 485938 484866 486174
rect 485102 485938 485134 486174
rect 484514 485854 485134 485938
rect 484514 485618 484546 485854
rect 484782 485618 484866 485854
rect 485102 485618 485134 485854
rect 484514 426174 485134 485618
rect 484514 425938 484546 426174
rect 484782 425938 484866 426174
rect 485102 425938 485134 426174
rect 484514 425854 485134 425938
rect 484514 425618 484546 425854
rect 484782 425618 484866 425854
rect 485102 425618 485134 425854
rect 484514 366174 485134 425618
rect 484514 365938 484546 366174
rect 484782 365938 484866 366174
rect 485102 365938 485134 366174
rect 484514 365854 485134 365938
rect 484514 365618 484546 365854
rect 484782 365618 484866 365854
rect 485102 365618 485134 365854
rect 484514 306174 485134 365618
rect 484514 305938 484546 306174
rect 484782 305938 484866 306174
rect 485102 305938 485134 306174
rect 484514 305854 485134 305938
rect 484514 305618 484546 305854
rect 484782 305618 484866 305854
rect 485102 305618 485134 305854
rect 484514 246174 485134 305618
rect 484514 245938 484546 246174
rect 484782 245938 484866 246174
rect 485102 245938 485134 246174
rect 484514 245854 485134 245938
rect 484514 245618 484546 245854
rect 484782 245618 484866 245854
rect 485102 245618 485134 245854
rect 484514 186174 485134 245618
rect 484514 185938 484546 186174
rect 484782 185938 484866 186174
rect 485102 185938 485134 186174
rect 484514 185854 485134 185938
rect 484514 185618 484546 185854
rect 484782 185618 484866 185854
rect 485102 185618 485134 185854
rect 484514 126174 485134 185618
rect 484514 125938 484546 126174
rect 484782 125938 484866 126174
rect 485102 125938 485134 126174
rect 484514 125854 485134 125938
rect 484514 125618 484546 125854
rect 484782 125618 484866 125854
rect 485102 125618 485134 125854
rect 484514 66174 485134 125618
rect 484514 65938 484546 66174
rect 484782 65938 484866 66174
rect 485102 65938 485134 66174
rect 484514 65854 485134 65938
rect 484514 65618 484546 65854
rect 484782 65618 484866 65854
rect 485102 65618 485134 65854
rect 484514 6174 485134 65618
rect 484514 5938 484546 6174
rect 484782 5938 484866 6174
rect 485102 5938 485134 6174
rect 484514 5854 485134 5938
rect 484514 5618 484546 5854
rect 484782 5618 484866 5854
rect 485102 5618 485134 5854
rect 484514 -2266 485134 5618
rect 484514 -2502 484546 -2266
rect 484782 -2502 484866 -2266
rect 485102 -2502 485134 -2266
rect 484514 -2586 485134 -2502
rect 484514 -2822 484546 -2586
rect 484782 -2822 484866 -2586
rect 485102 -2822 485134 -2586
rect 484514 -3814 485134 -2822
rect 488234 669894 488854 708122
rect 488234 669658 488266 669894
rect 488502 669658 488586 669894
rect 488822 669658 488854 669894
rect 488234 669574 488854 669658
rect 488234 669338 488266 669574
rect 488502 669338 488586 669574
rect 488822 669338 488854 669574
rect 488234 609894 488854 669338
rect 488234 609658 488266 609894
rect 488502 609658 488586 609894
rect 488822 609658 488854 609894
rect 488234 609574 488854 609658
rect 488234 609338 488266 609574
rect 488502 609338 488586 609574
rect 488822 609338 488854 609574
rect 488234 549894 488854 609338
rect 488234 549658 488266 549894
rect 488502 549658 488586 549894
rect 488822 549658 488854 549894
rect 488234 549574 488854 549658
rect 488234 549338 488266 549574
rect 488502 549338 488586 549574
rect 488822 549338 488854 549574
rect 488234 489894 488854 549338
rect 488234 489658 488266 489894
rect 488502 489658 488586 489894
rect 488822 489658 488854 489894
rect 488234 489574 488854 489658
rect 488234 489338 488266 489574
rect 488502 489338 488586 489574
rect 488822 489338 488854 489574
rect 488234 429894 488854 489338
rect 488234 429658 488266 429894
rect 488502 429658 488586 429894
rect 488822 429658 488854 429894
rect 488234 429574 488854 429658
rect 488234 429338 488266 429574
rect 488502 429338 488586 429574
rect 488822 429338 488854 429574
rect 488234 369894 488854 429338
rect 488234 369658 488266 369894
rect 488502 369658 488586 369894
rect 488822 369658 488854 369894
rect 488234 369574 488854 369658
rect 488234 369338 488266 369574
rect 488502 369338 488586 369574
rect 488822 369338 488854 369574
rect 488234 309894 488854 369338
rect 488234 309658 488266 309894
rect 488502 309658 488586 309894
rect 488822 309658 488854 309894
rect 488234 309574 488854 309658
rect 488234 309338 488266 309574
rect 488502 309338 488586 309574
rect 488822 309338 488854 309574
rect 488234 249894 488854 309338
rect 488234 249658 488266 249894
rect 488502 249658 488586 249894
rect 488822 249658 488854 249894
rect 488234 249574 488854 249658
rect 488234 249338 488266 249574
rect 488502 249338 488586 249574
rect 488822 249338 488854 249574
rect 488234 189894 488854 249338
rect 488234 189658 488266 189894
rect 488502 189658 488586 189894
rect 488822 189658 488854 189894
rect 488234 189574 488854 189658
rect 488234 189338 488266 189574
rect 488502 189338 488586 189574
rect 488822 189338 488854 189574
rect 488234 129894 488854 189338
rect 488234 129658 488266 129894
rect 488502 129658 488586 129894
rect 488822 129658 488854 129894
rect 488234 129574 488854 129658
rect 488234 129338 488266 129574
rect 488502 129338 488586 129574
rect 488822 129338 488854 129574
rect 488234 69894 488854 129338
rect 488234 69658 488266 69894
rect 488502 69658 488586 69894
rect 488822 69658 488854 69894
rect 488234 69574 488854 69658
rect 488234 69338 488266 69574
rect 488502 69338 488586 69574
rect 488822 69338 488854 69574
rect 488234 9894 488854 69338
rect 488234 9658 488266 9894
rect 488502 9658 488586 9894
rect 488822 9658 488854 9894
rect 488234 9574 488854 9658
rect 488234 9338 488266 9574
rect 488502 9338 488586 9574
rect 488822 9338 488854 9574
rect 488234 -4186 488854 9338
rect 488234 -4422 488266 -4186
rect 488502 -4422 488586 -4186
rect 488822 -4422 488854 -4186
rect 488234 -4506 488854 -4422
rect 488234 -4742 488266 -4506
rect 488502 -4742 488586 -4506
rect 488822 -4742 488854 -4506
rect 488234 -5734 488854 -4742
rect 491954 673614 492574 710042
rect 521954 711558 522574 711590
rect 521954 711322 521986 711558
rect 522222 711322 522306 711558
rect 522542 711322 522574 711558
rect 521954 711238 522574 711322
rect 521954 711002 521986 711238
rect 522222 711002 522306 711238
rect 522542 711002 522574 711238
rect 518234 709638 518854 709670
rect 518234 709402 518266 709638
rect 518502 709402 518586 709638
rect 518822 709402 518854 709638
rect 518234 709318 518854 709402
rect 518234 709082 518266 709318
rect 518502 709082 518586 709318
rect 518822 709082 518854 709318
rect 514514 707718 515134 707750
rect 514514 707482 514546 707718
rect 514782 707482 514866 707718
rect 515102 707482 515134 707718
rect 514514 707398 515134 707482
rect 514514 707162 514546 707398
rect 514782 707162 514866 707398
rect 515102 707162 515134 707398
rect 491954 673378 491986 673614
rect 492222 673378 492306 673614
rect 492542 673378 492574 673614
rect 491954 673294 492574 673378
rect 491954 673058 491986 673294
rect 492222 673058 492306 673294
rect 492542 673058 492574 673294
rect 491954 613614 492574 673058
rect 491954 613378 491986 613614
rect 492222 613378 492306 613614
rect 492542 613378 492574 613614
rect 491954 613294 492574 613378
rect 491954 613058 491986 613294
rect 492222 613058 492306 613294
rect 492542 613058 492574 613294
rect 491954 553614 492574 613058
rect 491954 553378 491986 553614
rect 492222 553378 492306 553614
rect 492542 553378 492574 553614
rect 491954 553294 492574 553378
rect 491954 553058 491986 553294
rect 492222 553058 492306 553294
rect 492542 553058 492574 553294
rect 491954 493614 492574 553058
rect 491954 493378 491986 493614
rect 492222 493378 492306 493614
rect 492542 493378 492574 493614
rect 491954 493294 492574 493378
rect 491954 493058 491986 493294
rect 492222 493058 492306 493294
rect 492542 493058 492574 493294
rect 491954 433614 492574 493058
rect 491954 433378 491986 433614
rect 492222 433378 492306 433614
rect 492542 433378 492574 433614
rect 491954 433294 492574 433378
rect 491954 433058 491986 433294
rect 492222 433058 492306 433294
rect 492542 433058 492574 433294
rect 491954 373614 492574 433058
rect 491954 373378 491986 373614
rect 492222 373378 492306 373614
rect 492542 373378 492574 373614
rect 491954 373294 492574 373378
rect 491954 373058 491986 373294
rect 492222 373058 492306 373294
rect 492542 373058 492574 373294
rect 491954 313614 492574 373058
rect 491954 313378 491986 313614
rect 492222 313378 492306 313614
rect 492542 313378 492574 313614
rect 491954 313294 492574 313378
rect 491954 313058 491986 313294
rect 492222 313058 492306 313294
rect 492542 313058 492574 313294
rect 491954 253614 492574 313058
rect 491954 253378 491986 253614
rect 492222 253378 492306 253614
rect 492542 253378 492574 253614
rect 491954 253294 492574 253378
rect 491954 253058 491986 253294
rect 492222 253058 492306 253294
rect 492542 253058 492574 253294
rect 491954 193614 492574 253058
rect 491954 193378 491986 193614
rect 492222 193378 492306 193614
rect 492542 193378 492574 193614
rect 491954 193294 492574 193378
rect 491954 193058 491986 193294
rect 492222 193058 492306 193294
rect 492542 193058 492574 193294
rect 491954 133614 492574 193058
rect 491954 133378 491986 133614
rect 492222 133378 492306 133614
rect 492542 133378 492574 133614
rect 491954 133294 492574 133378
rect 491954 133058 491986 133294
rect 492222 133058 492306 133294
rect 492542 133058 492574 133294
rect 491954 73614 492574 133058
rect 491954 73378 491986 73614
rect 492222 73378 492306 73614
rect 492542 73378 492574 73614
rect 491954 73294 492574 73378
rect 491954 73058 491986 73294
rect 492222 73058 492306 73294
rect 492542 73058 492574 73294
rect 491954 13614 492574 73058
rect 491954 13378 491986 13614
rect 492222 13378 492306 13614
rect 492542 13378 492574 13614
rect 491954 13294 492574 13378
rect 491954 13058 491986 13294
rect 492222 13058 492306 13294
rect 492542 13058 492574 13294
rect 461954 -7302 461986 -7066
rect 462222 -7302 462306 -7066
rect 462542 -7302 462574 -7066
rect 461954 -7386 462574 -7302
rect 461954 -7622 461986 -7386
rect 462222 -7622 462306 -7386
rect 462542 -7622 462574 -7386
rect 461954 -7654 462574 -7622
rect 491954 -6106 492574 13058
rect 510794 705798 511414 705830
rect 510794 705562 510826 705798
rect 511062 705562 511146 705798
rect 511382 705562 511414 705798
rect 510794 705478 511414 705562
rect 510794 705242 510826 705478
rect 511062 705242 511146 705478
rect 511382 705242 511414 705478
rect 510794 692454 511414 705242
rect 510794 692218 510826 692454
rect 511062 692218 511146 692454
rect 511382 692218 511414 692454
rect 510794 692134 511414 692218
rect 510794 691898 510826 692134
rect 511062 691898 511146 692134
rect 511382 691898 511414 692134
rect 510794 632454 511414 691898
rect 510794 632218 510826 632454
rect 511062 632218 511146 632454
rect 511382 632218 511414 632454
rect 510794 632134 511414 632218
rect 510794 631898 510826 632134
rect 511062 631898 511146 632134
rect 511382 631898 511414 632134
rect 510794 572454 511414 631898
rect 510794 572218 510826 572454
rect 511062 572218 511146 572454
rect 511382 572218 511414 572454
rect 510794 572134 511414 572218
rect 510794 571898 510826 572134
rect 511062 571898 511146 572134
rect 511382 571898 511414 572134
rect 510794 512454 511414 571898
rect 510794 512218 510826 512454
rect 511062 512218 511146 512454
rect 511382 512218 511414 512454
rect 510794 512134 511414 512218
rect 510794 511898 510826 512134
rect 511062 511898 511146 512134
rect 511382 511898 511414 512134
rect 510794 452454 511414 511898
rect 510794 452218 510826 452454
rect 511062 452218 511146 452454
rect 511382 452218 511414 452454
rect 510794 452134 511414 452218
rect 510794 451898 510826 452134
rect 511062 451898 511146 452134
rect 511382 451898 511414 452134
rect 510794 392454 511414 451898
rect 510794 392218 510826 392454
rect 511062 392218 511146 392454
rect 511382 392218 511414 392454
rect 510794 392134 511414 392218
rect 510794 391898 510826 392134
rect 511062 391898 511146 392134
rect 511382 391898 511414 392134
rect 510794 332454 511414 391898
rect 510794 332218 510826 332454
rect 511062 332218 511146 332454
rect 511382 332218 511414 332454
rect 510794 332134 511414 332218
rect 510794 331898 510826 332134
rect 511062 331898 511146 332134
rect 511382 331898 511414 332134
rect 510794 272454 511414 331898
rect 510794 272218 510826 272454
rect 511062 272218 511146 272454
rect 511382 272218 511414 272454
rect 510794 272134 511414 272218
rect 510794 271898 510826 272134
rect 511062 271898 511146 272134
rect 511382 271898 511414 272134
rect 510794 212454 511414 271898
rect 510794 212218 510826 212454
rect 511062 212218 511146 212454
rect 511382 212218 511414 212454
rect 510794 212134 511414 212218
rect 510794 211898 510826 212134
rect 511062 211898 511146 212134
rect 511382 211898 511414 212134
rect 510794 152454 511414 211898
rect 510794 152218 510826 152454
rect 511062 152218 511146 152454
rect 511382 152218 511414 152454
rect 510794 152134 511414 152218
rect 510794 151898 510826 152134
rect 511062 151898 511146 152134
rect 511382 151898 511414 152134
rect 510794 92454 511414 151898
rect 510794 92218 510826 92454
rect 511062 92218 511146 92454
rect 511382 92218 511414 92454
rect 510794 92134 511414 92218
rect 510794 91898 510826 92134
rect 511062 91898 511146 92134
rect 511382 91898 511414 92134
rect 510794 32454 511414 91898
rect 510794 32218 510826 32454
rect 511062 32218 511146 32454
rect 511382 32218 511414 32454
rect 510794 32134 511414 32218
rect 510794 31898 510826 32134
rect 511062 31898 511146 32134
rect 511382 31898 511414 32134
rect 510794 -1306 511414 31898
rect 510794 -1542 510826 -1306
rect 511062 -1542 511146 -1306
rect 511382 -1542 511414 -1306
rect 510794 -1626 511414 -1542
rect 510794 -1862 510826 -1626
rect 511062 -1862 511146 -1626
rect 511382 -1862 511414 -1626
rect 510794 -1894 511414 -1862
rect 514514 696174 515134 707162
rect 514514 695938 514546 696174
rect 514782 695938 514866 696174
rect 515102 695938 515134 696174
rect 514514 695854 515134 695938
rect 514514 695618 514546 695854
rect 514782 695618 514866 695854
rect 515102 695618 515134 695854
rect 514514 636174 515134 695618
rect 514514 635938 514546 636174
rect 514782 635938 514866 636174
rect 515102 635938 515134 636174
rect 514514 635854 515134 635938
rect 514514 635618 514546 635854
rect 514782 635618 514866 635854
rect 515102 635618 515134 635854
rect 514514 576174 515134 635618
rect 514514 575938 514546 576174
rect 514782 575938 514866 576174
rect 515102 575938 515134 576174
rect 514514 575854 515134 575938
rect 514514 575618 514546 575854
rect 514782 575618 514866 575854
rect 515102 575618 515134 575854
rect 514514 516174 515134 575618
rect 514514 515938 514546 516174
rect 514782 515938 514866 516174
rect 515102 515938 515134 516174
rect 514514 515854 515134 515938
rect 514514 515618 514546 515854
rect 514782 515618 514866 515854
rect 515102 515618 515134 515854
rect 514514 456174 515134 515618
rect 514514 455938 514546 456174
rect 514782 455938 514866 456174
rect 515102 455938 515134 456174
rect 514514 455854 515134 455938
rect 514514 455618 514546 455854
rect 514782 455618 514866 455854
rect 515102 455618 515134 455854
rect 514514 396174 515134 455618
rect 514514 395938 514546 396174
rect 514782 395938 514866 396174
rect 515102 395938 515134 396174
rect 514514 395854 515134 395938
rect 514514 395618 514546 395854
rect 514782 395618 514866 395854
rect 515102 395618 515134 395854
rect 514514 336174 515134 395618
rect 514514 335938 514546 336174
rect 514782 335938 514866 336174
rect 515102 335938 515134 336174
rect 514514 335854 515134 335938
rect 514514 335618 514546 335854
rect 514782 335618 514866 335854
rect 515102 335618 515134 335854
rect 514514 276174 515134 335618
rect 514514 275938 514546 276174
rect 514782 275938 514866 276174
rect 515102 275938 515134 276174
rect 514514 275854 515134 275938
rect 514514 275618 514546 275854
rect 514782 275618 514866 275854
rect 515102 275618 515134 275854
rect 514514 216174 515134 275618
rect 514514 215938 514546 216174
rect 514782 215938 514866 216174
rect 515102 215938 515134 216174
rect 514514 215854 515134 215938
rect 514514 215618 514546 215854
rect 514782 215618 514866 215854
rect 515102 215618 515134 215854
rect 514514 156174 515134 215618
rect 514514 155938 514546 156174
rect 514782 155938 514866 156174
rect 515102 155938 515134 156174
rect 514514 155854 515134 155938
rect 514514 155618 514546 155854
rect 514782 155618 514866 155854
rect 515102 155618 515134 155854
rect 514514 96174 515134 155618
rect 514514 95938 514546 96174
rect 514782 95938 514866 96174
rect 515102 95938 515134 96174
rect 514514 95854 515134 95938
rect 514514 95618 514546 95854
rect 514782 95618 514866 95854
rect 515102 95618 515134 95854
rect 514514 36174 515134 95618
rect 514514 35938 514546 36174
rect 514782 35938 514866 36174
rect 515102 35938 515134 36174
rect 514514 35854 515134 35938
rect 514514 35618 514546 35854
rect 514782 35618 514866 35854
rect 515102 35618 515134 35854
rect 514514 -3226 515134 35618
rect 514514 -3462 514546 -3226
rect 514782 -3462 514866 -3226
rect 515102 -3462 515134 -3226
rect 514514 -3546 515134 -3462
rect 514514 -3782 514546 -3546
rect 514782 -3782 514866 -3546
rect 515102 -3782 515134 -3546
rect 514514 -3814 515134 -3782
rect 518234 699894 518854 709082
rect 518234 699658 518266 699894
rect 518502 699658 518586 699894
rect 518822 699658 518854 699894
rect 518234 699574 518854 699658
rect 518234 699338 518266 699574
rect 518502 699338 518586 699574
rect 518822 699338 518854 699574
rect 518234 639894 518854 699338
rect 518234 639658 518266 639894
rect 518502 639658 518586 639894
rect 518822 639658 518854 639894
rect 518234 639574 518854 639658
rect 518234 639338 518266 639574
rect 518502 639338 518586 639574
rect 518822 639338 518854 639574
rect 518234 579894 518854 639338
rect 518234 579658 518266 579894
rect 518502 579658 518586 579894
rect 518822 579658 518854 579894
rect 518234 579574 518854 579658
rect 518234 579338 518266 579574
rect 518502 579338 518586 579574
rect 518822 579338 518854 579574
rect 518234 519894 518854 579338
rect 518234 519658 518266 519894
rect 518502 519658 518586 519894
rect 518822 519658 518854 519894
rect 518234 519574 518854 519658
rect 518234 519338 518266 519574
rect 518502 519338 518586 519574
rect 518822 519338 518854 519574
rect 518234 459894 518854 519338
rect 518234 459658 518266 459894
rect 518502 459658 518586 459894
rect 518822 459658 518854 459894
rect 518234 459574 518854 459658
rect 518234 459338 518266 459574
rect 518502 459338 518586 459574
rect 518822 459338 518854 459574
rect 518234 399894 518854 459338
rect 518234 399658 518266 399894
rect 518502 399658 518586 399894
rect 518822 399658 518854 399894
rect 518234 399574 518854 399658
rect 518234 399338 518266 399574
rect 518502 399338 518586 399574
rect 518822 399338 518854 399574
rect 518234 339894 518854 399338
rect 518234 339658 518266 339894
rect 518502 339658 518586 339894
rect 518822 339658 518854 339894
rect 518234 339574 518854 339658
rect 518234 339338 518266 339574
rect 518502 339338 518586 339574
rect 518822 339338 518854 339574
rect 518234 279894 518854 339338
rect 518234 279658 518266 279894
rect 518502 279658 518586 279894
rect 518822 279658 518854 279894
rect 518234 279574 518854 279658
rect 518234 279338 518266 279574
rect 518502 279338 518586 279574
rect 518822 279338 518854 279574
rect 518234 219894 518854 279338
rect 518234 219658 518266 219894
rect 518502 219658 518586 219894
rect 518822 219658 518854 219894
rect 518234 219574 518854 219658
rect 518234 219338 518266 219574
rect 518502 219338 518586 219574
rect 518822 219338 518854 219574
rect 518234 159894 518854 219338
rect 518234 159658 518266 159894
rect 518502 159658 518586 159894
rect 518822 159658 518854 159894
rect 518234 159574 518854 159658
rect 518234 159338 518266 159574
rect 518502 159338 518586 159574
rect 518822 159338 518854 159574
rect 518234 99894 518854 159338
rect 518234 99658 518266 99894
rect 518502 99658 518586 99894
rect 518822 99658 518854 99894
rect 518234 99574 518854 99658
rect 518234 99338 518266 99574
rect 518502 99338 518586 99574
rect 518822 99338 518854 99574
rect 518234 39894 518854 99338
rect 518234 39658 518266 39894
rect 518502 39658 518586 39894
rect 518822 39658 518854 39894
rect 518234 39574 518854 39658
rect 518234 39338 518266 39574
rect 518502 39338 518586 39574
rect 518822 39338 518854 39574
rect 518234 -5146 518854 39338
rect 518234 -5382 518266 -5146
rect 518502 -5382 518586 -5146
rect 518822 -5382 518854 -5146
rect 518234 -5466 518854 -5382
rect 518234 -5702 518266 -5466
rect 518502 -5702 518586 -5466
rect 518822 -5702 518854 -5466
rect 518234 -5734 518854 -5702
rect 521954 643614 522574 711002
rect 551954 710598 552574 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 551954 710362 551986 710598
rect 552222 710362 552306 710598
rect 552542 710362 552574 710598
rect 551954 710278 552574 710362
rect 551954 710042 551986 710278
rect 552222 710042 552306 710278
rect 552542 710042 552574 710278
rect 548234 708678 548854 709670
rect 548234 708442 548266 708678
rect 548502 708442 548586 708678
rect 548822 708442 548854 708678
rect 548234 708358 548854 708442
rect 548234 708122 548266 708358
rect 548502 708122 548586 708358
rect 548822 708122 548854 708358
rect 544514 706758 545134 707750
rect 544514 706522 544546 706758
rect 544782 706522 544866 706758
rect 545102 706522 545134 706758
rect 544514 706438 545134 706522
rect 544514 706202 544546 706438
rect 544782 706202 544866 706438
rect 545102 706202 545134 706438
rect 521954 643378 521986 643614
rect 522222 643378 522306 643614
rect 522542 643378 522574 643614
rect 521954 643294 522574 643378
rect 521954 643058 521986 643294
rect 522222 643058 522306 643294
rect 522542 643058 522574 643294
rect 521954 583614 522574 643058
rect 521954 583378 521986 583614
rect 522222 583378 522306 583614
rect 522542 583378 522574 583614
rect 521954 583294 522574 583378
rect 521954 583058 521986 583294
rect 522222 583058 522306 583294
rect 522542 583058 522574 583294
rect 521954 523614 522574 583058
rect 521954 523378 521986 523614
rect 522222 523378 522306 523614
rect 522542 523378 522574 523614
rect 521954 523294 522574 523378
rect 521954 523058 521986 523294
rect 522222 523058 522306 523294
rect 522542 523058 522574 523294
rect 521954 463614 522574 523058
rect 521954 463378 521986 463614
rect 522222 463378 522306 463614
rect 522542 463378 522574 463614
rect 521954 463294 522574 463378
rect 521954 463058 521986 463294
rect 522222 463058 522306 463294
rect 522542 463058 522574 463294
rect 521954 403614 522574 463058
rect 521954 403378 521986 403614
rect 522222 403378 522306 403614
rect 522542 403378 522574 403614
rect 521954 403294 522574 403378
rect 521954 403058 521986 403294
rect 522222 403058 522306 403294
rect 522542 403058 522574 403294
rect 521954 343614 522574 403058
rect 521954 343378 521986 343614
rect 522222 343378 522306 343614
rect 522542 343378 522574 343614
rect 521954 343294 522574 343378
rect 521954 343058 521986 343294
rect 522222 343058 522306 343294
rect 522542 343058 522574 343294
rect 521954 283614 522574 343058
rect 521954 283378 521986 283614
rect 522222 283378 522306 283614
rect 522542 283378 522574 283614
rect 521954 283294 522574 283378
rect 521954 283058 521986 283294
rect 522222 283058 522306 283294
rect 522542 283058 522574 283294
rect 521954 223614 522574 283058
rect 521954 223378 521986 223614
rect 522222 223378 522306 223614
rect 522542 223378 522574 223614
rect 521954 223294 522574 223378
rect 521954 223058 521986 223294
rect 522222 223058 522306 223294
rect 522542 223058 522574 223294
rect 521954 163614 522574 223058
rect 521954 163378 521986 163614
rect 522222 163378 522306 163614
rect 522542 163378 522574 163614
rect 521954 163294 522574 163378
rect 521954 163058 521986 163294
rect 522222 163058 522306 163294
rect 522542 163058 522574 163294
rect 521954 103614 522574 163058
rect 521954 103378 521986 103614
rect 522222 103378 522306 103614
rect 522542 103378 522574 103614
rect 521954 103294 522574 103378
rect 521954 103058 521986 103294
rect 522222 103058 522306 103294
rect 522542 103058 522574 103294
rect 521954 43614 522574 103058
rect 521954 43378 521986 43614
rect 522222 43378 522306 43614
rect 522542 43378 522574 43614
rect 521954 43294 522574 43378
rect 521954 43058 521986 43294
rect 522222 43058 522306 43294
rect 522542 43058 522574 43294
rect 491954 -6342 491986 -6106
rect 492222 -6342 492306 -6106
rect 492542 -6342 492574 -6106
rect 491954 -6426 492574 -6342
rect 491954 -6662 491986 -6426
rect 492222 -6662 492306 -6426
rect 492542 -6662 492574 -6426
rect 491954 -7654 492574 -6662
rect 521954 -7066 522574 43058
rect 540794 704838 541414 705830
rect 540794 704602 540826 704838
rect 541062 704602 541146 704838
rect 541382 704602 541414 704838
rect 540794 704518 541414 704602
rect 540794 704282 540826 704518
rect 541062 704282 541146 704518
rect 541382 704282 541414 704518
rect 540794 662454 541414 704282
rect 540794 662218 540826 662454
rect 541062 662218 541146 662454
rect 541382 662218 541414 662454
rect 540794 662134 541414 662218
rect 540794 661898 540826 662134
rect 541062 661898 541146 662134
rect 541382 661898 541414 662134
rect 540794 602454 541414 661898
rect 540794 602218 540826 602454
rect 541062 602218 541146 602454
rect 541382 602218 541414 602454
rect 540794 602134 541414 602218
rect 540794 601898 540826 602134
rect 541062 601898 541146 602134
rect 541382 601898 541414 602134
rect 540794 542454 541414 601898
rect 540794 542218 540826 542454
rect 541062 542218 541146 542454
rect 541382 542218 541414 542454
rect 540794 542134 541414 542218
rect 540794 541898 540826 542134
rect 541062 541898 541146 542134
rect 541382 541898 541414 542134
rect 540794 482454 541414 541898
rect 540794 482218 540826 482454
rect 541062 482218 541146 482454
rect 541382 482218 541414 482454
rect 540794 482134 541414 482218
rect 540794 481898 540826 482134
rect 541062 481898 541146 482134
rect 541382 481898 541414 482134
rect 540794 422454 541414 481898
rect 540794 422218 540826 422454
rect 541062 422218 541146 422454
rect 541382 422218 541414 422454
rect 540794 422134 541414 422218
rect 540794 421898 540826 422134
rect 541062 421898 541146 422134
rect 541382 421898 541414 422134
rect 540794 362454 541414 421898
rect 540794 362218 540826 362454
rect 541062 362218 541146 362454
rect 541382 362218 541414 362454
rect 540794 362134 541414 362218
rect 540794 361898 540826 362134
rect 541062 361898 541146 362134
rect 541382 361898 541414 362134
rect 540794 302454 541414 361898
rect 540794 302218 540826 302454
rect 541062 302218 541146 302454
rect 541382 302218 541414 302454
rect 540794 302134 541414 302218
rect 540794 301898 540826 302134
rect 541062 301898 541146 302134
rect 541382 301898 541414 302134
rect 540794 242454 541414 301898
rect 540794 242218 540826 242454
rect 541062 242218 541146 242454
rect 541382 242218 541414 242454
rect 540794 242134 541414 242218
rect 540794 241898 540826 242134
rect 541062 241898 541146 242134
rect 541382 241898 541414 242134
rect 540794 182454 541414 241898
rect 540794 182218 540826 182454
rect 541062 182218 541146 182454
rect 541382 182218 541414 182454
rect 540794 182134 541414 182218
rect 540794 181898 540826 182134
rect 541062 181898 541146 182134
rect 541382 181898 541414 182134
rect 540794 122454 541414 181898
rect 540794 122218 540826 122454
rect 541062 122218 541146 122454
rect 541382 122218 541414 122454
rect 540794 122134 541414 122218
rect 540794 121898 540826 122134
rect 541062 121898 541146 122134
rect 541382 121898 541414 122134
rect 540794 62454 541414 121898
rect 540794 62218 540826 62454
rect 541062 62218 541146 62454
rect 541382 62218 541414 62454
rect 540794 62134 541414 62218
rect 540794 61898 540826 62134
rect 541062 61898 541146 62134
rect 541382 61898 541414 62134
rect 540794 2454 541414 61898
rect 540794 2218 540826 2454
rect 541062 2218 541146 2454
rect 541382 2218 541414 2454
rect 540794 2134 541414 2218
rect 540794 1898 540826 2134
rect 541062 1898 541146 2134
rect 541382 1898 541414 2134
rect 540794 -346 541414 1898
rect 540794 -582 540826 -346
rect 541062 -582 541146 -346
rect 541382 -582 541414 -346
rect 540794 -666 541414 -582
rect 540794 -902 540826 -666
rect 541062 -902 541146 -666
rect 541382 -902 541414 -666
rect 540794 -1894 541414 -902
rect 544514 666174 545134 706202
rect 544514 665938 544546 666174
rect 544782 665938 544866 666174
rect 545102 665938 545134 666174
rect 544514 665854 545134 665938
rect 544514 665618 544546 665854
rect 544782 665618 544866 665854
rect 545102 665618 545134 665854
rect 544514 606174 545134 665618
rect 544514 605938 544546 606174
rect 544782 605938 544866 606174
rect 545102 605938 545134 606174
rect 544514 605854 545134 605938
rect 544514 605618 544546 605854
rect 544782 605618 544866 605854
rect 545102 605618 545134 605854
rect 544514 546174 545134 605618
rect 544514 545938 544546 546174
rect 544782 545938 544866 546174
rect 545102 545938 545134 546174
rect 544514 545854 545134 545938
rect 544514 545618 544546 545854
rect 544782 545618 544866 545854
rect 545102 545618 545134 545854
rect 544514 486174 545134 545618
rect 544514 485938 544546 486174
rect 544782 485938 544866 486174
rect 545102 485938 545134 486174
rect 544514 485854 545134 485938
rect 544514 485618 544546 485854
rect 544782 485618 544866 485854
rect 545102 485618 545134 485854
rect 544514 426174 545134 485618
rect 544514 425938 544546 426174
rect 544782 425938 544866 426174
rect 545102 425938 545134 426174
rect 544514 425854 545134 425938
rect 544514 425618 544546 425854
rect 544782 425618 544866 425854
rect 545102 425618 545134 425854
rect 544514 366174 545134 425618
rect 544514 365938 544546 366174
rect 544782 365938 544866 366174
rect 545102 365938 545134 366174
rect 544514 365854 545134 365938
rect 544514 365618 544546 365854
rect 544782 365618 544866 365854
rect 545102 365618 545134 365854
rect 544514 306174 545134 365618
rect 544514 305938 544546 306174
rect 544782 305938 544866 306174
rect 545102 305938 545134 306174
rect 544514 305854 545134 305938
rect 544514 305618 544546 305854
rect 544782 305618 544866 305854
rect 545102 305618 545134 305854
rect 544514 246174 545134 305618
rect 544514 245938 544546 246174
rect 544782 245938 544866 246174
rect 545102 245938 545134 246174
rect 544514 245854 545134 245938
rect 544514 245618 544546 245854
rect 544782 245618 544866 245854
rect 545102 245618 545134 245854
rect 544514 186174 545134 245618
rect 544514 185938 544546 186174
rect 544782 185938 544866 186174
rect 545102 185938 545134 186174
rect 544514 185854 545134 185938
rect 544514 185618 544546 185854
rect 544782 185618 544866 185854
rect 545102 185618 545134 185854
rect 544514 126174 545134 185618
rect 544514 125938 544546 126174
rect 544782 125938 544866 126174
rect 545102 125938 545134 126174
rect 544514 125854 545134 125938
rect 544514 125618 544546 125854
rect 544782 125618 544866 125854
rect 545102 125618 545134 125854
rect 544514 66174 545134 125618
rect 544514 65938 544546 66174
rect 544782 65938 544866 66174
rect 545102 65938 545134 66174
rect 544514 65854 545134 65938
rect 544514 65618 544546 65854
rect 544782 65618 544866 65854
rect 545102 65618 545134 65854
rect 544514 6174 545134 65618
rect 544514 5938 544546 6174
rect 544782 5938 544866 6174
rect 545102 5938 545134 6174
rect 544514 5854 545134 5938
rect 544514 5618 544546 5854
rect 544782 5618 544866 5854
rect 545102 5618 545134 5854
rect 544514 -2266 545134 5618
rect 544514 -2502 544546 -2266
rect 544782 -2502 544866 -2266
rect 545102 -2502 545134 -2266
rect 544514 -2586 545134 -2502
rect 544514 -2822 544546 -2586
rect 544782 -2822 544866 -2586
rect 545102 -2822 545134 -2586
rect 544514 -3814 545134 -2822
rect 548234 669894 548854 708122
rect 548234 669658 548266 669894
rect 548502 669658 548586 669894
rect 548822 669658 548854 669894
rect 548234 669574 548854 669658
rect 548234 669338 548266 669574
rect 548502 669338 548586 669574
rect 548822 669338 548854 669574
rect 548234 609894 548854 669338
rect 548234 609658 548266 609894
rect 548502 609658 548586 609894
rect 548822 609658 548854 609894
rect 548234 609574 548854 609658
rect 548234 609338 548266 609574
rect 548502 609338 548586 609574
rect 548822 609338 548854 609574
rect 548234 549894 548854 609338
rect 548234 549658 548266 549894
rect 548502 549658 548586 549894
rect 548822 549658 548854 549894
rect 548234 549574 548854 549658
rect 548234 549338 548266 549574
rect 548502 549338 548586 549574
rect 548822 549338 548854 549574
rect 548234 489894 548854 549338
rect 548234 489658 548266 489894
rect 548502 489658 548586 489894
rect 548822 489658 548854 489894
rect 548234 489574 548854 489658
rect 548234 489338 548266 489574
rect 548502 489338 548586 489574
rect 548822 489338 548854 489574
rect 548234 429894 548854 489338
rect 548234 429658 548266 429894
rect 548502 429658 548586 429894
rect 548822 429658 548854 429894
rect 548234 429574 548854 429658
rect 548234 429338 548266 429574
rect 548502 429338 548586 429574
rect 548822 429338 548854 429574
rect 548234 369894 548854 429338
rect 548234 369658 548266 369894
rect 548502 369658 548586 369894
rect 548822 369658 548854 369894
rect 548234 369574 548854 369658
rect 548234 369338 548266 369574
rect 548502 369338 548586 369574
rect 548822 369338 548854 369574
rect 548234 309894 548854 369338
rect 548234 309658 548266 309894
rect 548502 309658 548586 309894
rect 548822 309658 548854 309894
rect 548234 309574 548854 309658
rect 548234 309338 548266 309574
rect 548502 309338 548586 309574
rect 548822 309338 548854 309574
rect 548234 249894 548854 309338
rect 548234 249658 548266 249894
rect 548502 249658 548586 249894
rect 548822 249658 548854 249894
rect 548234 249574 548854 249658
rect 548234 249338 548266 249574
rect 548502 249338 548586 249574
rect 548822 249338 548854 249574
rect 548234 189894 548854 249338
rect 548234 189658 548266 189894
rect 548502 189658 548586 189894
rect 548822 189658 548854 189894
rect 548234 189574 548854 189658
rect 548234 189338 548266 189574
rect 548502 189338 548586 189574
rect 548822 189338 548854 189574
rect 548234 129894 548854 189338
rect 548234 129658 548266 129894
rect 548502 129658 548586 129894
rect 548822 129658 548854 129894
rect 548234 129574 548854 129658
rect 548234 129338 548266 129574
rect 548502 129338 548586 129574
rect 548822 129338 548854 129574
rect 548234 69894 548854 129338
rect 548234 69658 548266 69894
rect 548502 69658 548586 69894
rect 548822 69658 548854 69894
rect 548234 69574 548854 69658
rect 548234 69338 548266 69574
rect 548502 69338 548586 69574
rect 548822 69338 548854 69574
rect 548234 9894 548854 69338
rect 548234 9658 548266 9894
rect 548502 9658 548586 9894
rect 548822 9658 548854 9894
rect 548234 9574 548854 9658
rect 548234 9338 548266 9574
rect 548502 9338 548586 9574
rect 548822 9338 548854 9574
rect 548234 -4186 548854 9338
rect 548234 -4422 548266 -4186
rect 548502 -4422 548586 -4186
rect 548822 -4422 548854 -4186
rect 548234 -4506 548854 -4422
rect 548234 -4742 548266 -4506
rect 548502 -4742 548586 -4506
rect 548822 -4742 548854 -4506
rect 548234 -5734 548854 -4742
rect 551954 673614 552574 710042
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 578234 709638 578854 709670
rect 578234 709402 578266 709638
rect 578502 709402 578586 709638
rect 578822 709402 578854 709638
rect 578234 709318 578854 709402
rect 578234 709082 578266 709318
rect 578502 709082 578586 709318
rect 578822 709082 578854 709318
rect 574514 707718 575134 707750
rect 574514 707482 574546 707718
rect 574782 707482 574866 707718
rect 575102 707482 575134 707718
rect 574514 707398 575134 707482
rect 574514 707162 574546 707398
rect 574782 707162 574866 707398
rect 575102 707162 575134 707398
rect 551954 673378 551986 673614
rect 552222 673378 552306 673614
rect 552542 673378 552574 673614
rect 551954 673294 552574 673378
rect 551954 673058 551986 673294
rect 552222 673058 552306 673294
rect 552542 673058 552574 673294
rect 551954 613614 552574 673058
rect 551954 613378 551986 613614
rect 552222 613378 552306 613614
rect 552542 613378 552574 613614
rect 551954 613294 552574 613378
rect 551954 613058 551986 613294
rect 552222 613058 552306 613294
rect 552542 613058 552574 613294
rect 551954 553614 552574 613058
rect 551954 553378 551986 553614
rect 552222 553378 552306 553614
rect 552542 553378 552574 553614
rect 551954 553294 552574 553378
rect 551954 553058 551986 553294
rect 552222 553058 552306 553294
rect 552542 553058 552574 553294
rect 551954 493614 552574 553058
rect 551954 493378 551986 493614
rect 552222 493378 552306 493614
rect 552542 493378 552574 493614
rect 551954 493294 552574 493378
rect 551954 493058 551986 493294
rect 552222 493058 552306 493294
rect 552542 493058 552574 493294
rect 551954 433614 552574 493058
rect 551954 433378 551986 433614
rect 552222 433378 552306 433614
rect 552542 433378 552574 433614
rect 551954 433294 552574 433378
rect 551954 433058 551986 433294
rect 552222 433058 552306 433294
rect 552542 433058 552574 433294
rect 551954 373614 552574 433058
rect 551954 373378 551986 373614
rect 552222 373378 552306 373614
rect 552542 373378 552574 373614
rect 551954 373294 552574 373378
rect 551954 373058 551986 373294
rect 552222 373058 552306 373294
rect 552542 373058 552574 373294
rect 551954 313614 552574 373058
rect 551954 313378 551986 313614
rect 552222 313378 552306 313614
rect 552542 313378 552574 313614
rect 551954 313294 552574 313378
rect 551954 313058 551986 313294
rect 552222 313058 552306 313294
rect 552542 313058 552574 313294
rect 551954 253614 552574 313058
rect 551954 253378 551986 253614
rect 552222 253378 552306 253614
rect 552542 253378 552574 253614
rect 551954 253294 552574 253378
rect 551954 253058 551986 253294
rect 552222 253058 552306 253294
rect 552542 253058 552574 253294
rect 551954 193614 552574 253058
rect 551954 193378 551986 193614
rect 552222 193378 552306 193614
rect 552542 193378 552574 193614
rect 551954 193294 552574 193378
rect 551954 193058 551986 193294
rect 552222 193058 552306 193294
rect 552542 193058 552574 193294
rect 551954 133614 552574 193058
rect 551954 133378 551986 133614
rect 552222 133378 552306 133614
rect 552542 133378 552574 133614
rect 551954 133294 552574 133378
rect 551954 133058 551986 133294
rect 552222 133058 552306 133294
rect 552542 133058 552574 133294
rect 551954 73614 552574 133058
rect 551954 73378 551986 73614
rect 552222 73378 552306 73614
rect 552542 73378 552574 73614
rect 551954 73294 552574 73378
rect 551954 73058 551986 73294
rect 552222 73058 552306 73294
rect 552542 73058 552574 73294
rect 551954 13614 552574 73058
rect 551954 13378 551986 13614
rect 552222 13378 552306 13614
rect 552542 13378 552574 13614
rect 551954 13294 552574 13378
rect 551954 13058 551986 13294
rect 552222 13058 552306 13294
rect 552542 13058 552574 13294
rect 521954 -7302 521986 -7066
rect 522222 -7302 522306 -7066
rect 522542 -7302 522574 -7066
rect 521954 -7386 522574 -7302
rect 521954 -7622 521986 -7386
rect 522222 -7622 522306 -7386
rect 522542 -7622 522574 -7386
rect 521954 -7654 522574 -7622
rect 551954 -6106 552574 13058
rect 570794 705798 571414 705830
rect 570794 705562 570826 705798
rect 571062 705562 571146 705798
rect 571382 705562 571414 705798
rect 570794 705478 571414 705562
rect 570794 705242 570826 705478
rect 571062 705242 571146 705478
rect 571382 705242 571414 705478
rect 570794 692454 571414 705242
rect 570794 692218 570826 692454
rect 571062 692218 571146 692454
rect 571382 692218 571414 692454
rect 570794 692134 571414 692218
rect 570794 691898 570826 692134
rect 571062 691898 571146 692134
rect 571382 691898 571414 692134
rect 570794 632454 571414 691898
rect 570794 632218 570826 632454
rect 571062 632218 571146 632454
rect 571382 632218 571414 632454
rect 570794 632134 571414 632218
rect 570794 631898 570826 632134
rect 571062 631898 571146 632134
rect 571382 631898 571414 632134
rect 570794 572454 571414 631898
rect 570794 572218 570826 572454
rect 571062 572218 571146 572454
rect 571382 572218 571414 572454
rect 570794 572134 571414 572218
rect 570794 571898 570826 572134
rect 571062 571898 571146 572134
rect 571382 571898 571414 572134
rect 570794 512454 571414 571898
rect 570794 512218 570826 512454
rect 571062 512218 571146 512454
rect 571382 512218 571414 512454
rect 570794 512134 571414 512218
rect 570794 511898 570826 512134
rect 571062 511898 571146 512134
rect 571382 511898 571414 512134
rect 570794 452454 571414 511898
rect 570794 452218 570826 452454
rect 571062 452218 571146 452454
rect 571382 452218 571414 452454
rect 570794 452134 571414 452218
rect 570794 451898 570826 452134
rect 571062 451898 571146 452134
rect 571382 451898 571414 452134
rect 570794 392454 571414 451898
rect 570794 392218 570826 392454
rect 571062 392218 571146 392454
rect 571382 392218 571414 392454
rect 570794 392134 571414 392218
rect 570794 391898 570826 392134
rect 571062 391898 571146 392134
rect 571382 391898 571414 392134
rect 570794 332454 571414 391898
rect 570794 332218 570826 332454
rect 571062 332218 571146 332454
rect 571382 332218 571414 332454
rect 570794 332134 571414 332218
rect 570794 331898 570826 332134
rect 571062 331898 571146 332134
rect 571382 331898 571414 332134
rect 570794 272454 571414 331898
rect 570794 272218 570826 272454
rect 571062 272218 571146 272454
rect 571382 272218 571414 272454
rect 570794 272134 571414 272218
rect 570794 271898 570826 272134
rect 571062 271898 571146 272134
rect 571382 271898 571414 272134
rect 570794 212454 571414 271898
rect 570794 212218 570826 212454
rect 571062 212218 571146 212454
rect 571382 212218 571414 212454
rect 570794 212134 571414 212218
rect 570794 211898 570826 212134
rect 571062 211898 571146 212134
rect 571382 211898 571414 212134
rect 570794 152454 571414 211898
rect 570794 152218 570826 152454
rect 571062 152218 571146 152454
rect 571382 152218 571414 152454
rect 570794 152134 571414 152218
rect 570794 151898 570826 152134
rect 571062 151898 571146 152134
rect 571382 151898 571414 152134
rect 570794 92454 571414 151898
rect 570794 92218 570826 92454
rect 571062 92218 571146 92454
rect 571382 92218 571414 92454
rect 570794 92134 571414 92218
rect 570794 91898 570826 92134
rect 571062 91898 571146 92134
rect 571382 91898 571414 92134
rect 570794 32454 571414 91898
rect 570794 32218 570826 32454
rect 571062 32218 571146 32454
rect 571382 32218 571414 32454
rect 570794 32134 571414 32218
rect 570794 31898 570826 32134
rect 571062 31898 571146 32134
rect 571382 31898 571414 32134
rect 570794 -1306 571414 31898
rect 570794 -1542 570826 -1306
rect 571062 -1542 571146 -1306
rect 571382 -1542 571414 -1306
rect 570794 -1626 571414 -1542
rect 570794 -1862 570826 -1626
rect 571062 -1862 571146 -1626
rect 571382 -1862 571414 -1626
rect 570794 -1894 571414 -1862
rect 574514 696174 575134 707162
rect 574514 695938 574546 696174
rect 574782 695938 574866 696174
rect 575102 695938 575134 696174
rect 574514 695854 575134 695938
rect 574514 695618 574546 695854
rect 574782 695618 574866 695854
rect 575102 695618 575134 695854
rect 574514 636174 575134 695618
rect 574514 635938 574546 636174
rect 574782 635938 574866 636174
rect 575102 635938 575134 636174
rect 574514 635854 575134 635938
rect 574514 635618 574546 635854
rect 574782 635618 574866 635854
rect 575102 635618 575134 635854
rect 574514 576174 575134 635618
rect 574514 575938 574546 576174
rect 574782 575938 574866 576174
rect 575102 575938 575134 576174
rect 574514 575854 575134 575938
rect 574514 575618 574546 575854
rect 574782 575618 574866 575854
rect 575102 575618 575134 575854
rect 574514 516174 575134 575618
rect 574514 515938 574546 516174
rect 574782 515938 574866 516174
rect 575102 515938 575134 516174
rect 574514 515854 575134 515938
rect 574514 515618 574546 515854
rect 574782 515618 574866 515854
rect 575102 515618 575134 515854
rect 574514 456174 575134 515618
rect 574514 455938 574546 456174
rect 574782 455938 574866 456174
rect 575102 455938 575134 456174
rect 574514 455854 575134 455938
rect 574514 455618 574546 455854
rect 574782 455618 574866 455854
rect 575102 455618 575134 455854
rect 574514 396174 575134 455618
rect 574514 395938 574546 396174
rect 574782 395938 574866 396174
rect 575102 395938 575134 396174
rect 574514 395854 575134 395938
rect 574514 395618 574546 395854
rect 574782 395618 574866 395854
rect 575102 395618 575134 395854
rect 574514 336174 575134 395618
rect 574514 335938 574546 336174
rect 574782 335938 574866 336174
rect 575102 335938 575134 336174
rect 574514 335854 575134 335938
rect 574514 335618 574546 335854
rect 574782 335618 574866 335854
rect 575102 335618 575134 335854
rect 574514 276174 575134 335618
rect 574514 275938 574546 276174
rect 574782 275938 574866 276174
rect 575102 275938 575134 276174
rect 574514 275854 575134 275938
rect 574514 275618 574546 275854
rect 574782 275618 574866 275854
rect 575102 275618 575134 275854
rect 574514 216174 575134 275618
rect 574514 215938 574546 216174
rect 574782 215938 574866 216174
rect 575102 215938 575134 216174
rect 574514 215854 575134 215938
rect 574514 215618 574546 215854
rect 574782 215618 574866 215854
rect 575102 215618 575134 215854
rect 574514 156174 575134 215618
rect 574514 155938 574546 156174
rect 574782 155938 574866 156174
rect 575102 155938 575134 156174
rect 574514 155854 575134 155938
rect 574514 155618 574546 155854
rect 574782 155618 574866 155854
rect 575102 155618 575134 155854
rect 574514 96174 575134 155618
rect 574514 95938 574546 96174
rect 574782 95938 574866 96174
rect 575102 95938 575134 96174
rect 574514 95854 575134 95938
rect 574514 95618 574546 95854
rect 574782 95618 574866 95854
rect 575102 95618 575134 95854
rect 574514 36174 575134 95618
rect 574514 35938 574546 36174
rect 574782 35938 574866 36174
rect 575102 35938 575134 36174
rect 574514 35854 575134 35938
rect 574514 35618 574546 35854
rect 574782 35618 574866 35854
rect 575102 35618 575134 35854
rect 574514 -3226 575134 35618
rect 574514 -3462 574546 -3226
rect 574782 -3462 574866 -3226
rect 575102 -3462 575134 -3226
rect 574514 -3546 575134 -3462
rect 574514 -3782 574546 -3546
rect 574782 -3782 574866 -3546
rect 575102 -3782 575134 -3546
rect 574514 -3814 575134 -3782
rect 578234 699894 578854 709082
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 578234 699658 578266 699894
rect 578502 699658 578586 699894
rect 578822 699658 578854 699894
rect 578234 699574 578854 699658
rect 578234 699338 578266 699574
rect 578502 699338 578586 699574
rect 578822 699338 578854 699574
rect 578234 639894 578854 699338
rect 578234 639658 578266 639894
rect 578502 639658 578586 639894
rect 578822 639658 578854 639894
rect 578234 639574 578854 639658
rect 578234 639338 578266 639574
rect 578502 639338 578586 639574
rect 578822 639338 578854 639574
rect 578234 579894 578854 639338
rect 578234 579658 578266 579894
rect 578502 579658 578586 579894
rect 578822 579658 578854 579894
rect 578234 579574 578854 579658
rect 578234 579338 578266 579574
rect 578502 579338 578586 579574
rect 578822 579338 578854 579574
rect 578234 519894 578854 579338
rect 578234 519658 578266 519894
rect 578502 519658 578586 519894
rect 578822 519658 578854 519894
rect 578234 519574 578854 519658
rect 578234 519338 578266 519574
rect 578502 519338 578586 519574
rect 578822 519338 578854 519574
rect 578234 459894 578854 519338
rect 578234 459658 578266 459894
rect 578502 459658 578586 459894
rect 578822 459658 578854 459894
rect 578234 459574 578854 459658
rect 578234 459338 578266 459574
rect 578502 459338 578586 459574
rect 578822 459338 578854 459574
rect 578234 399894 578854 459338
rect 578234 399658 578266 399894
rect 578502 399658 578586 399894
rect 578822 399658 578854 399894
rect 578234 399574 578854 399658
rect 578234 399338 578266 399574
rect 578502 399338 578586 399574
rect 578822 399338 578854 399574
rect 578234 339894 578854 399338
rect 578234 339658 578266 339894
rect 578502 339658 578586 339894
rect 578822 339658 578854 339894
rect 578234 339574 578854 339658
rect 578234 339338 578266 339574
rect 578502 339338 578586 339574
rect 578822 339338 578854 339574
rect 578234 279894 578854 339338
rect 578234 279658 578266 279894
rect 578502 279658 578586 279894
rect 578822 279658 578854 279894
rect 578234 279574 578854 279658
rect 578234 279338 578266 279574
rect 578502 279338 578586 279574
rect 578822 279338 578854 279574
rect 578234 219894 578854 279338
rect 578234 219658 578266 219894
rect 578502 219658 578586 219894
rect 578822 219658 578854 219894
rect 578234 219574 578854 219658
rect 578234 219338 578266 219574
rect 578502 219338 578586 219574
rect 578822 219338 578854 219574
rect 578234 159894 578854 219338
rect 578234 159658 578266 159894
rect 578502 159658 578586 159894
rect 578822 159658 578854 159894
rect 578234 159574 578854 159658
rect 578234 159338 578266 159574
rect 578502 159338 578586 159574
rect 578822 159338 578854 159574
rect 578234 99894 578854 159338
rect 578234 99658 578266 99894
rect 578502 99658 578586 99894
rect 578822 99658 578854 99894
rect 578234 99574 578854 99658
rect 578234 99338 578266 99574
rect 578502 99338 578586 99574
rect 578822 99338 578854 99574
rect 578234 39894 578854 99338
rect 578234 39658 578266 39894
rect 578502 39658 578586 39894
rect 578822 39658 578854 39894
rect 578234 39574 578854 39658
rect 578234 39338 578266 39574
rect 578502 39338 578586 39574
rect 578822 39338 578854 39574
rect 578234 -5146 578854 39338
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 662454 585930 704282
rect 585310 662218 585342 662454
rect 585578 662218 585662 662454
rect 585898 662218 585930 662454
rect 585310 662134 585930 662218
rect 585310 661898 585342 662134
rect 585578 661898 585662 662134
rect 585898 661898 585930 662134
rect 585310 602454 585930 661898
rect 585310 602218 585342 602454
rect 585578 602218 585662 602454
rect 585898 602218 585930 602454
rect 585310 602134 585930 602218
rect 585310 601898 585342 602134
rect 585578 601898 585662 602134
rect 585898 601898 585930 602134
rect 585310 542454 585930 601898
rect 585310 542218 585342 542454
rect 585578 542218 585662 542454
rect 585898 542218 585930 542454
rect 585310 542134 585930 542218
rect 585310 541898 585342 542134
rect 585578 541898 585662 542134
rect 585898 541898 585930 542134
rect 585310 482454 585930 541898
rect 585310 482218 585342 482454
rect 585578 482218 585662 482454
rect 585898 482218 585930 482454
rect 585310 482134 585930 482218
rect 585310 481898 585342 482134
rect 585578 481898 585662 482134
rect 585898 481898 585930 482134
rect 585310 422454 585930 481898
rect 585310 422218 585342 422454
rect 585578 422218 585662 422454
rect 585898 422218 585930 422454
rect 585310 422134 585930 422218
rect 585310 421898 585342 422134
rect 585578 421898 585662 422134
rect 585898 421898 585930 422134
rect 585310 362454 585930 421898
rect 585310 362218 585342 362454
rect 585578 362218 585662 362454
rect 585898 362218 585930 362454
rect 585310 362134 585930 362218
rect 585310 361898 585342 362134
rect 585578 361898 585662 362134
rect 585898 361898 585930 362134
rect 585310 302454 585930 361898
rect 585310 302218 585342 302454
rect 585578 302218 585662 302454
rect 585898 302218 585930 302454
rect 585310 302134 585930 302218
rect 585310 301898 585342 302134
rect 585578 301898 585662 302134
rect 585898 301898 585930 302134
rect 585310 242454 585930 301898
rect 585310 242218 585342 242454
rect 585578 242218 585662 242454
rect 585898 242218 585930 242454
rect 585310 242134 585930 242218
rect 585310 241898 585342 242134
rect 585578 241898 585662 242134
rect 585898 241898 585930 242134
rect 585310 182454 585930 241898
rect 585310 182218 585342 182454
rect 585578 182218 585662 182454
rect 585898 182218 585930 182454
rect 585310 182134 585930 182218
rect 585310 181898 585342 182134
rect 585578 181898 585662 182134
rect 585898 181898 585930 182134
rect 585310 122454 585930 181898
rect 585310 122218 585342 122454
rect 585578 122218 585662 122454
rect 585898 122218 585930 122454
rect 585310 122134 585930 122218
rect 585310 121898 585342 122134
rect 585578 121898 585662 122134
rect 585898 121898 585930 122134
rect 585310 62454 585930 121898
rect 585310 62218 585342 62454
rect 585578 62218 585662 62454
rect 585898 62218 585930 62454
rect 585310 62134 585930 62218
rect 585310 61898 585342 62134
rect 585578 61898 585662 62134
rect 585898 61898 585930 62134
rect 585310 2454 585930 61898
rect 585310 2218 585342 2454
rect 585578 2218 585662 2454
rect 585898 2218 585930 2454
rect 585310 2134 585930 2218
rect 585310 1898 585342 2134
rect 585578 1898 585662 2134
rect 585898 1898 585930 2134
rect 585310 -346 585930 1898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 692454 586890 705242
rect 586270 692218 586302 692454
rect 586538 692218 586622 692454
rect 586858 692218 586890 692454
rect 586270 692134 586890 692218
rect 586270 691898 586302 692134
rect 586538 691898 586622 692134
rect 586858 691898 586890 692134
rect 586270 632454 586890 691898
rect 586270 632218 586302 632454
rect 586538 632218 586622 632454
rect 586858 632218 586890 632454
rect 586270 632134 586890 632218
rect 586270 631898 586302 632134
rect 586538 631898 586622 632134
rect 586858 631898 586890 632134
rect 586270 572454 586890 631898
rect 586270 572218 586302 572454
rect 586538 572218 586622 572454
rect 586858 572218 586890 572454
rect 586270 572134 586890 572218
rect 586270 571898 586302 572134
rect 586538 571898 586622 572134
rect 586858 571898 586890 572134
rect 586270 512454 586890 571898
rect 586270 512218 586302 512454
rect 586538 512218 586622 512454
rect 586858 512218 586890 512454
rect 586270 512134 586890 512218
rect 586270 511898 586302 512134
rect 586538 511898 586622 512134
rect 586858 511898 586890 512134
rect 586270 452454 586890 511898
rect 586270 452218 586302 452454
rect 586538 452218 586622 452454
rect 586858 452218 586890 452454
rect 586270 452134 586890 452218
rect 586270 451898 586302 452134
rect 586538 451898 586622 452134
rect 586858 451898 586890 452134
rect 586270 392454 586890 451898
rect 586270 392218 586302 392454
rect 586538 392218 586622 392454
rect 586858 392218 586890 392454
rect 586270 392134 586890 392218
rect 586270 391898 586302 392134
rect 586538 391898 586622 392134
rect 586858 391898 586890 392134
rect 586270 332454 586890 391898
rect 586270 332218 586302 332454
rect 586538 332218 586622 332454
rect 586858 332218 586890 332454
rect 586270 332134 586890 332218
rect 586270 331898 586302 332134
rect 586538 331898 586622 332134
rect 586858 331898 586890 332134
rect 586270 272454 586890 331898
rect 586270 272218 586302 272454
rect 586538 272218 586622 272454
rect 586858 272218 586890 272454
rect 586270 272134 586890 272218
rect 586270 271898 586302 272134
rect 586538 271898 586622 272134
rect 586858 271898 586890 272134
rect 586270 212454 586890 271898
rect 586270 212218 586302 212454
rect 586538 212218 586622 212454
rect 586858 212218 586890 212454
rect 586270 212134 586890 212218
rect 586270 211898 586302 212134
rect 586538 211898 586622 212134
rect 586858 211898 586890 212134
rect 586270 152454 586890 211898
rect 586270 152218 586302 152454
rect 586538 152218 586622 152454
rect 586858 152218 586890 152454
rect 586270 152134 586890 152218
rect 586270 151898 586302 152134
rect 586538 151898 586622 152134
rect 586858 151898 586890 152134
rect 586270 92454 586890 151898
rect 586270 92218 586302 92454
rect 586538 92218 586622 92454
rect 586858 92218 586890 92454
rect 586270 92134 586890 92218
rect 586270 91898 586302 92134
rect 586538 91898 586622 92134
rect 586858 91898 586890 92134
rect 586270 32454 586890 91898
rect 586270 32218 586302 32454
rect 586538 32218 586622 32454
rect 586858 32218 586890 32454
rect 586270 32134 586890 32218
rect 586270 31898 586302 32134
rect 586538 31898 586622 32134
rect 586858 31898 586890 32134
rect 586270 -1306 586890 31898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 666174 587850 706202
rect 587230 665938 587262 666174
rect 587498 665938 587582 666174
rect 587818 665938 587850 666174
rect 587230 665854 587850 665938
rect 587230 665618 587262 665854
rect 587498 665618 587582 665854
rect 587818 665618 587850 665854
rect 587230 606174 587850 665618
rect 587230 605938 587262 606174
rect 587498 605938 587582 606174
rect 587818 605938 587850 606174
rect 587230 605854 587850 605938
rect 587230 605618 587262 605854
rect 587498 605618 587582 605854
rect 587818 605618 587850 605854
rect 587230 546174 587850 605618
rect 587230 545938 587262 546174
rect 587498 545938 587582 546174
rect 587818 545938 587850 546174
rect 587230 545854 587850 545938
rect 587230 545618 587262 545854
rect 587498 545618 587582 545854
rect 587818 545618 587850 545854
rect 587230 486174 587850 545618
rect 587230 485938 587262 486174
rect 587498 485938 587582 486174
rect 587818 485938 587850 486174
rect 587230 485854 587850 485938
rect 587230 485618 587262 485854
rect 587498 485618 587582 485854
rect 587818 485618 587850 485854
rect 587230 426174 587850 485618
rect 587230 425938 587262 426174
rect 587498 425938 587582 426174
rect 587818 425938 587850 426174
rect 587230 425854 587850 425938
rect 587230 425618 587262 425854
rect 587498 425618 587582 425854
rect 587818 425618 587850 425854
rect 587230 366174 587850 425618
rect 587230 365938 587262 366174
rect 587498 365938 587582 366174
rect 587818 365938 587850 366174
rect 587230 365854 587850 365938
rect 587230 365618 587262 365854
rect 587498 365618 587582 365854
rect 587818 365618 587850 365854
rect 587230 306174 587850 365618
rect 587230 305938 587262 306174
rect 587498 305938 587582 306174
rect 587818 305938 587850 306174
rect 587230 305854 587850 305938
rect 587230 305618 587262 305854
rect 587498 305618 587582 305854
rect 587818 305618 587850 305854
rect 587230 246174 587850 305618
rect 587230 245938 587262 246174
rect 587498 245938 587582 246174
rect 587818 245938 587850 246174
rect 587230 245854 587850 245938
rect 587230 245618 587262 245854
rect 587498 245618 587582 245854
rect 587818 245618 587850 245854
rect 587230 186174 587850 245618
rect 587230 185938 587262 186174
rect 587498 185938 587582 186174
rect 587818 185938 587850 186174
rect 587230 185854 587850 185938
rect 587230 185618 587262 185854
rect 587498 185618 587582 185854
rect 587818 185618 587850 185854
rect 587230 126174 587850 185618
rect 587230 125938 587262 126174
rect 587498 125938 587582 126174
rect 587818 125938 587850 126174
rect 587230 125854 587850 125938
rect 587230 125618 587262 125854
rect 587498 125618 587582 125854
rect 587818 125618 587850 125854
rect 587230 66174 587850 125618
rect 587230 65938 587262 66174
rect 587498 65938 587582 66174
rect 587818 65938 587850 66174
rect 587230 65854 587850 65938
rect 587230 65618 587262 65854
rect 587498 65618 587582 65854
rect 587818 65618 587850 65854
rect 587230 6174 587850 65618
rect 587230 5938 587262 6174
rect 587498 5938 587582 6174
rect 587818 5938 587850 6174
rect 587230 5854 587850 5938
rect 587230 5618 587262 5854
rect 587498 5618 587582 5854
rect 587818 5618 587850 5854
rect 587230 -2266 587850 5618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 696174 588810 707162
rect 588190 695938 588222 696174
rect 588458 695938 588542 696174
rect 588778 695938 588810 696174
rect 588190 695854 588810 695938
rect 588190 695618 588222 695854
rect 588458 695618 588542 695854
rect 588778 695618 588810 695854
rect 588190 636174 588810 695618
rect 588190 635938 588222 636174
rect 588458 635938 588542 636174
rect 588778 635938 588810 636174
rect 588190 635854 588810 635938
rect 588190 635618 588222 635854
rect 588458 635618 588542 635854
rect 588778 635618 588810 635854
rect 588190 576174 588810 635618
rect 588190 575938 588222 576174
rect 588458 575938 588542 576174
rect 588778 575938 588810 576174
rect 588190 575854 588810 575938
rect 588190 575618 588222 575854
rect 588458 575618 588542 575854
rect 588778 575618 588810 575854
rect 588190 516174 588810 575618
rect 588190 515938 588222 516174
rect 588458 515938 588542 516174
rect 588778 515938 588810 516174
rect 588190 515854 588810 515938
rect 588190 515618 588222 515854
rect 588458 515618 588542 515854
rect 588778 515618 588810 515854
rect 588190 456174 588810 515618
rect 588190 455938 588222 456174
rect 588458 455938 588542 456174
rect 588778 455938 588810 456174
rect 588190 455854 588810 455938
rect 588190 455618 588222 455854
rect 588458 455618 588542 455854
rect 588778 455618 588810 455854
rect 588190 396174 588810 455618
rect 588190 395938 588222 396174
rect 588458 395938 588542 396174
rect 588778 395938 588810 396174
rect 588190 395854 588810 395938
rect 588190 395618 588222 395854
rect 588458 395618 588542 395854
rect 588778 395618 588810 395854
rect 588190 336174 588810 395618
rect 588190 335938 588222 336174
rect 588458 335938 588542 336174
rect 588778 335938 588810 336174
rect 588190 335854 588810 335938
rect 588190 335618 588222 335854
rect 588458 335618 588542 335854
rect 588778 335618 588810 335854
rect 588190 276174 588810 335618
rect 588190 275938 588222 276174
rect 588458 275938 588542 276174
rect 588778 275938 588810 276174
rect 588190 275854 588810 275938
rect 588190 275618 588222 275854
rect 588458 275618 588542 275854
rect 588778 275618 588810 275854
rect 588190 216174 588810 275618
rect 588190 215938 588222 216174
rect 588458 215938 588542 216174
rect 588778 215938 588810 216174
rect 588190 215854 588810 215938
rect 588190 215618 588222 215854
rect 588458 215618 588542 215854
rect 588778 215618 588810 215854
rect 588190 156174 588810 215618
rect 588190 155938 588222 156174
rect 588458 155938 588542 156174
rect 588778 155938 588810 156174
rect 588190 155854 588810 155938
rect 588190 155618 588222 155854
rect 588458 155618 588542 155854
rect 588778 155618 588810 155854
rect 588190 96174 588810 155618
rect 588190 95938 588222 96174
rect 588458 95938 588542 96174
rect 588778 95938 588810 96174
rect 588190 95854 588810 95938
rect 588190 95618 588222 95854
rect 588458 95618 588542 95854
rect 588778 95618 588810 95854
rect 588190 36174 588810 95618
rect 588190 35938 588222 36174
rect 588458 35938 588542 36174
rect 588778 35938 588810 36174
rect 588190 35854 588810 35938
rect 588190 35618 588222 35854
rect 588458 35618 588542 35854
rect 588778 35618 588810 35854
rect 588190 -3226 588810 35618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669894 589770 708122
rect 589150 669658 589182 669894
rect 589418 669658 589502 669894
rect 589738 669658 589770 669894
rect 589150 669574 589770 669658
rect 589150 669338 589182 669574
rect 589418 669338 589502 669574
rect 589738 669338 589770 669574
rect 589150 609894 589770 669338
rect 589150 609658 589182 609894
rect 589418 609658 589502 609894
rect 589738 609658 589770 609894
rect 589150 609574 589770 609658
rect 589150 609338 589182 609574
rect 589418 609338 589502 609574
rect 589738 609338 589770 609574
rect 589150 549894 589770 609338
rect 589150 549658 589182 549894
rect 589418 549658 589502 549894
rect 589738 549658 589770 549894
rect 589150 549574 589770 549658
rect 589150 549338 589182 549574
rect 589418 549338 589502 549574
rect 589738 549338 589770 549574
rect 589150 489894 589770 549338
rect 589150 489658 589182 489894
rect 589418 489658 589502 489894
rect 589738 489658 589770 489894
rect 589150 489574 589770 489658
rect 589150 489338 589182 489574
rect 589418 489338 589502 489574
rect 589738 489338 589770 489574
rect 589150 429894 589770 489338
rect 589150 429658 589182 429894
rect 589418 429658 589502 429894
rect 589738 429658 589770 429894
rect 589150 429574 589770 429658
rect 589150 429338 589182 429574
rect 589418 429338 589502 429574
rect 589738 429338 589770 429574
rect 589150 369894 589770 429338
rect 589150 369658 589182 369894
rect 589418 369658 589502 369894
rect 589738 369658 589770 369894
rect 589150 369574 589770 369658
rect 589150 369338 589182 369574
rect 589418 369338 589502 369574
rect 589738 369338 589770 369574
rect 589150 309894 589770 369338
rect 589150 309658 589182 309894
rect 589418 309658 589502 309894
rect 589738 309658 589770 309894
rect 589150 309574 589770 309658
rect 589150 309338 589182 309574
rect 589418 309338 589502 309574
rect 589738 309338 589770 309574
rect 589150 249894 589770 309338
rect 589150 249658 589182 249894
rect 589418 249658 589502 249894
rect 589738 249658 589770 249894
rect 589150 249574 589770 249658
rect 589150 249338 589182 249574
rect 589418 249338 589502 249574
rect 589738 249338 589770 249574
rect 589150 189894 589770 249338
rect 589150 189658 589182 189894
rect 589418 189658 589502 189894
rect 589738 189658 589770 189894
rect 589150 189574 589770 189658
rect 589150 189338 589182 189574
rect 589418 189338 589502 189574
rect 589738 189338 589770 189574
rect 589150 129894 589770 189338
rect 589150 129658 589182 129894
rect 589418 129658 589502 129894
rect 589738 129658 589770 129894
rect 589150 129574 589770 129658
rect 589150 129338 589182 129574
rect 589418 129338 589502 129574
rect 589738 129338 589770 129574
rect 589150 69894 589770 129338
rect 589150 69658 589182 69894
rect 589418 69658 589502 69894
rect 589738 69658 589770 69894
rect 589150 69574 589770 69658
rect 589150 69338 589182 69574
rect 589418 69338 589502 69574
rect 589738 69338 589770 69574
rect 589150 9894 589770 69338
rect 589150 9658 589182 9894
rect 589418 9658 589502 9894
rect 589738 9658 589770 9894
rect 589150 9574 589770 9658
rect 589150 9338 589182 9574
rect 589418 9338 589502 9574
rect 589738 9338 589770 9574
rect 589150 -4186 589770 9338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 699894 590730 709082
rect 590110 699658 590142 699894
rect 590378 699658 590462 699894
rect 590698 699658 590730 699894
rect 590110 699574 590730 699658
rect 590110 699338 590142 699574
rect 590378 699338 590462 699574
rect 590698 699338 590730 699574
rect 590110 639894 590730 699338
rect 590110 639658 590142 639894
rect 590378 639658 590462 639894
rect 590698 639658 590730 639894
rect 590110 639574 590730 639658
rect 590110 639338 590142 639574
rect 590378 639338 590462 639574
rect 590698 639338 590730 639574
rect 590110 579894 590730 639338
rect 590110 579658 590142 579894
rect 590378 579658 590462 579894
rect 590698 579658 590730 579894
rect 590110 579574 590730 579658
rect 590110 579338 590142 579574
rect 590378 579338 590462 579574
rect 590698 579338 590730 579574
rect 590110 519894 590730 579338
rect 590110 519658 590142 519894
rect 590378 519658 590462 519894
rect 590698 519658 590730 519894
rect 590110 519574 590730 519658
rect 590110 519338 590142 519574
rect 590378 519338 590462 519574
rect 590698 519338 590730 519574
rect 590110 459894 590730 519338
rect 590110 459658 590142 459894
rect 590378 459658 590462 459894
rect 590698 459658 590730 459894
rect 590110 459574 590730 459658
rect 590110 459338 590142 459574
rect 590378 459338 590462 459574
rect 590698 459338 590730 459574
rect 590110 399894 590730 459338
rect 590110 399658 590142 399894
rect 590378 399658 590462 399894
rect 590698 399658 590730 399894
rect 590110 399574 590730 399658
rect 590110 399338 590142 399574
rect 590378 399338 590462 399574
rect 590698 399338 590730 399574
rect 590110 339894 590730 399338
rect 590110 339658 590142 339894
rect 590378 339658 590462 339894
rect 590698 339658 590730 339894
rect 590110 339574 590730 339658
rect 590110 339338 590142 339574
rect 590378 339338 590462 339574
rect 590698 339338 590730 339574
rect 590110 279894 590730 339338
rect 590110 279658 590142 279894
rect 590378 279658 590462 279894
rect 590698 279658 590730 279894
rect 590110 279574 590730 279658
rect 590110 279338 590142 279574
rect 590378 279338 590462 279574
rect 590698 279338 590730 279574
rect 590110 219894 590730 279338
rect 590110 219658 590142 219894
rect 590378 219658 590462 219894
rect 590698 219658 590730 219894
rect 590110 219574 590730 219658
rect 590110 219338 590142 219574
rect 590378 219338 590462 219574
rect 590698 219338 590730 219574
rect 590110 159894 590730 219338
rect 590110 159658 590142 159894
rect 590378 159658 590462 159894
rect 590698 159658 590730 159894
rect 590110 159574 590730 159658
rect 590110 159338 590142 159574
rect 590378 159338 590462 159574
rect 590698 159338 590730 159574
rect 590110 99894 590730 159338
rect 590110 99658 590142 99894
rect 590378 99658 590462 99894
rect 590698 99658 590730 99894
rect 590110 99574 590730 99658
rect 590110 99338 590142 99574
rect 590378 99338 590462 99574
rect 590698 99338 590730 99574
rect 590110 39894 590730 99338
rect 590110 39658 590142 39894
rect 590378 39658 590462 39894
rect 590698 39658 590730 39894
rect 590110 39574 590730 39658
rect 590110 39338 590142 39574
rect 590378 39338 590462 39574
rect 590698 39338 590730 39574
rect 578234 -5382 578266 -5146
rect 578502 -5382 578586 -5146
rect 578822 -5382 578854 -5146
rect 578234 -5466 578854 -5382
rect 578234 -5702 578266 -5466
rect 578502 -5702 578586 -5466
rect 578822 -5702 578854 -5466
rect 578234 -5734 578854 -5702
rect 590110 -5146 590730 39338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673614 591690 710042
rect 591070 673378 591102 673614
rect 591338 673378 591422 673614
rect 591658 673378 591690 673614
rect 591070 673294 591690 673378
rect 591070 673058 591102 673294
rect 591338 673058 591422 673294
rect 591658 673058 591690 673294
rect 591070 613614 591690 673058
rect 591070 613378 591102 613614
rect 591338 613378 591422 613614
rect 591658 613378 591690 613614
rect 591070 613294 591690 613378
rect 591070 613058 591102 613294
rect 591338 613058 591422 613294
rect 591658 613058 591690 613294
rect 591070 553614 591690 613058
rect 591070 553378 591102 553614
rect 591338 553378 591422 553614
rect 591658 553378 591690 553614
rect 591070 553294 591690 553378
rect 591070 553058 591102 553294
rect 591338 553058 591422 553294
rect 591658 553058 591690 553294
rect 591070 493614 591690 553058
rect 591070 493378 591102 493614
rect 591338 493378 591422 493614
rect 591658 493378 591690 493614
rect 591070 493294 591690 493378
rect 591070 493058 591102 493294
rect 591338 493058 591422 493294
rect 591658 493058 591690 493294
rect 591070 433614 591690 493058
rect 591070 433378 591102 433614
rect 591338 433378 591422 433614
rect 591658 433378 591690 433614
rect 591070 433294 591690 433378
rect 591070 433058 591102 433294
rect 591338 433058 591422 433294
rect 591658 433058 591690 433294
rect 591070 373614 591690 433058
rect 591070 373378 591102 373614
rect 591338 373378 591422 373614
rect 591658 373378 591690 373614
rect 591070 373294 591690 373378
rect 591070 373058 591102 373294
rect 591338 373058 591422 373294
rect 591658 373058 591690 373294
rect 591070 313614 591690 373058
rect 591070 313378 591102 313614
rect 591338 313378 591422 313614
rect 591658 313378 591690 313614
rect 591070 313294 591690 313378
rect 591070 313058 591102 313294
rect 591338 313058 591422 313294
rect 591658 313058 591690 313294
rect 591070 253614 591690 313058
rect 591070 253378 591102 253614
rect 591338 253378 591422 253614
rect 591658 253378 591690 253614
rect 591070 253294 591690 253378
rect 591070 253058 591102 253294
rect 591338 253058 591422 253294
rect 591658 253058 591690 253294
rect 591070 193614 591690 253058
rect 591070 193378 591102 193614
rect 591338 193378 591422 193614
rect 591658 193378 591690 193614
rect 591070 193294 591690 193378
rect 591070 193058 591102 193294
rect 591338 193058 591422 193294
rect 591658 193058 591690 193294
rect 591070 133614 591690 193058
rect 591070 133378 591102 133614
rect 591338 133378 591422 133614
rect 591658 133378 591690 133614
rect 591070 133294 591690 133378
rect 591070 133058 591102 133294
rect 591338 133058 591422 133294
rect 591658 133058 591690 133294
rect 591070 73614 591690 133058
rect 591070 73378 591102 73614
rect 591338 73378 591422 73614
rect 591658 73378 591690 73614
rect 591070 73294 591690 73378
rect 591070 73058 591102 73294
rect 591338 73058 591422 73294
rect 591658 73058 591690 73294
rect 591070 13614 591690 73058
rect 591070 13378 591102 13614
rect 591338 13378 591422 13614
rect 591658 13378 591690 13614
rect 591070 13294 591690 13378
rect 591070 13058 591102 13294
rect 591338 13058 591422 13294
rect 591658 13058 591690 13294
rect 551954 -6342 551986 -6106
rect 552222 -6342 552306 -6106
rect 552542 -6342 552574 -6106
rect 551954 -6426 552574 -6342
rect 551954 -6662 551986 -6426
rect 552222 -6662 552306 -6426
rect 552542 -6662 552574 -6426
rect 551954 -7654 552574 -6662
rect 591070 -6106 591690 13058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 643614 592650 711002
rect 592030 643378 592062 643614
rect 592298 643378 592382 643614
rect 592618 643378 592650 643614
rect 592030 643294 592650 643378
rect 592030 643058 592062 643294
rect 592298 643058 592382 643294
rect 592618 643058 592650 643294
rect 592030 583614 592650 643058
rect 592030 583378 592062 583614
rect 592298 583378 592382 583614
rect 592618 583378 592650 583614
rect 592030 583294 592650 583378
rect 592030 583058 592062 583294
rect 592298 583058 592382 583294
rect 592618 583058 592650 583294
rect 592030 523614 592650 583058
rect 592030 523378 592062 523614
rect 592298 523378 592382 523614
rect 592618 523378 592650 523614
rect 592030 523294 592650 523378
rect 592030 523058 592062 523294
rect 592298 523058 592382 523294
rect 592618 523058 592650 523294
rect 592030 463614 592650 523058
rect 592030 463378 592062 463614
rect 592298 463378 592382 463614
rect 592618 463378 592650 463614
rect 592030 463294 592650 463378
rect 592030 463058 592062 463294
rect 592298 463058 592382 463294
rect 592618 463058 592650 463294
rect 592030 403614 592650 463058
rect 592030 403378 592062 403614
rect 592298 403378 592382 403614
rect 592618 403378 592650 403614
rect 592030 403294 592650 403378
rect 592030 403058 592062 403294
rect 592298 403058 592382 403294
rect 592618 403058 592650 403294
rect 592030 343614 592650 403058
rect 592030 343378 592062 343614
rect 592298 343378 592382 343614
rect 592618 343378 592650 343614
rect 592030 343294 592650 343378
rect 592030 343058 592062 343294
rect 592298 343058 592382 343294
rect 592618 343058 592650 343294
rect 592030 283614 592650 343058
rect 592030 283378 592062 283614
rect 592298 283378 592382 283614
rect 592618 283378 592650 283614
rect 592030 283294 592650 283378
rect 592030 283058 592062 283294
rect 592298 283058 592382 283294
rect 592618 283058 592650 283294
rect 592030 223614 592650 283058
rect 592030 223378 592062 223614
rect 592298 223378 592382 223614
rect 592618 223378 592650 223614
rect 592030 223294 592650 223378
rect 592030 223058 592062 223294
rect 592298 223058 592382 223294
rect 592618 223058 592650 223294
rect 592030 163614 592650 223058
rect 592030 163378 592062 163614
rect 592298 163378 592382 163614
rect 592618 163378 592650 163614
rect 592030 163294 592650 163378
rect 592030 163058 592062 163294
rect 592298 163058 592382 163294
rect 592618 163058 592650 163294
rect 592030 103614 592650 163058
rect 592030 103378 592062 103614
rect 592298 103378 592382 103614
rect 592618 103378 592650 103614
rect 592030 103294 592650 103378
rect 592030 103058 592062 103294
rect 592298 103058 592382 103294
rect 592618 103058 592650 103294
rect 592030 43614 592650 103058
rect 592030 43378 592062 43614
rect 592298 43378 592382 43614
rect 592618 43378 592650 43614
rect 592030 43294 592650 43378
rect 592030 43058 592062 43294
rect 592298 43058 592382 43294
rect 592618 43058 592650 43294
rect 592030 -7066 592650 43058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 643378 -8458 643614
rect -8374 643378 -8138 643614
rect -8694 643058 -8458 643294
rect -8374 643058 -8138 643294
rect -8694 583378 -8458 583614
rect -8374 583378 -8138 583614
rect -8694 583058 -8458 583294
rect -8374 583058 -8138 583294
rect -8694 523378 -8458 523614
rect -8374 523378 -8138 523614
rect -8694 523058 -8458 523294
rect -8374 523058 -8138 523294
rect -8694 463378 -8458 463614
rect -8374 463378 -8138 463614
rect -8694 463058 -8458 463294
rect -8374 463058 -8138 463294
rect -8694 403378 -8458 403614
rect -8374 403378 -8138 403614
rect -8694 403058 -8458 403294
rect -8374 403058 -8138 403294
rect -8694 343378 -8458 343614
rect -8374 343378 -8138 343614
rect -8694 343058 -8458 343294
rect -8374 343058 -8138 343294
rect -8694 283378 -8458 283614
rect -8374 283378 -8138 283614
rect -8694 283058 -8458 283294
rect -8374 283058 -8138 283294
rect -8694 223378 -8458 223614
rect -8374 223378 -8138 223614
rect -8694 223058 -8458 223294
rect -8374 223058 -8138 223294
rect -8694 163378 -8458 163614
rect -8374 163378 -8138 163614
rect -8694 163058 -8458 163294
rect -8374 163058 -8138 163294
rect -8694 103378 -8458 103614
rect -8374 103378 -8138 103614
rect -8694 103058 -8458 103294
rect -8374 103058 -8138 103294
rect -8694 43378 -8458 43614
rect -8374 43378 -8138 43614
rect -8694 43058 -8458 43294
rect -8374 43058 -8138 43294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 11986 710362 12222 710598
rect 12306 710362 12542 710598
rect 11986 710042 12222 710278
rect 12306 710042 12542 710278
rect -7734 673378 -7498 673614
rect -7414 673378 -7178 673614
rect -7734 673058 -7498 673294
rect -7414 673058 -7178 673294
rect -7734 613378 -7498 613614
rect -7414 613378 -7178 613614
rect -7734 613058 -7498 613294
rect -7414 613058 -7178 613294
rect -7734 553378 -7498 553614
rect -7414 553378 -7178 553614
rect -7734 553058 -7498 553294
rect -7414 553058 -7178 553294
rect -7734 493378 -7498 493614
rect -7414 493378 -7178 493614
rect -7734 493058 -7498 493294
rect -7414 493058 -7178 493294
rect -7734 433378 -7498 433614
rect -7414 433378 -7178 433614
rect -7734 433058 -7498 433294
rect -7414 433058 -7178 433294
rect -7734 373378 -7498 373614
rect -7414 373378 -7178 373614
rect -7734 373058 -7498 373294
rect -7414 373058 -7178 373294
rect -7734 313378 -7498 313614
rect -7414 313378 -7178 313614
rect -7734 313058 -7498 313294
rect -7414 313058 -7178 313294
rect -7734 253378 -7498 253614
rect -7414 253378 -7178 253614
rect -7734 253058 -7498 253294
rect -7414 253058 -7178 253294
rect -7734 193378 -7498 193614
rect -7414 193378 -7178 193614
rect -7734 193058 -7498 193294
rect -7414 193058 -7178 193294
rect -7734 133378 -7498 133614
rect -7414 133378 -7178 133614
rect -7734 133058 -7498 133294
rect -7414 133058 -7178 133294
rect -7734 73378 -7498 73614
rect -7414 73378 -7178 73614
rect -7734 73058 -7498 73294
rect -7414 73058 -7178 73294
rect -7734 13378 -7498 13614
rect -7414 13378 -7178 13614
rect -7734 13058 -7498 13294
rect -7414 13058 -7178 13294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 699658 -6538 699894
rect -6454 699658 -6218 699894
rect -6774 699338 -6538 699574
rect -6454 699338 -6218 699574
rect -6774 639658 -6538 639894
rect -6454 639658 -6218 639894
rect -6774 639338 -6538 639574
rect -6454 639338 -6218 639574
rect -6774 579658 -6538 579894
rect -6454 579658 -6218 579894
rect -6774 579338 -6538 579574
rect -6454 579338 -6218 579574
rect -6774 519658 -6538 519894
rect -6454 519658 -6218 519894
rect -6774 519338 -6538 519574
rect -6454 519338 -6218 519574
rect -6774 459658 -6538 459894
rect -6454 459658 -6218 459894
rect -6774 459338 -6538 459574
rect -6454 459338 -6218 459574
rect -6774 399658 -6538 399894
rect -6454 399658 -6218 399894
rect -6774 399338 -6538 399574
rect -6454 399338 -6218 399574
rect -6774 339658 -6538 339894
rect -6454 339658 -6218 339894
rect -6774 339338 -6538 339574
rect -6454 339338 -6218 339574
rect -6774 279658 -6538 279894
rect -6454 279658 -6218 279894
rect -6774 279338 -6538 279574
rect -6454 279338 -6218 279574
rect -6774 219658 -6538 219894
rect -6454 219658 -6218 219894
rect -6774 219338 -6538 219574
rect -6454 219338 -6218 219574
rect -6774 159658 -6538 159894
rect -6454 159658 -6218 159894
rect -6774 159338 -6538 159574
rect -6454 159338 -6218 159574
rect -6774 99658 -6538 99894
rect -6454 99658 -6218 99894
rect -6774 99338 -6538 99574
rect -6454 99338 -6218 99574
rect -6774 39658 -6538 39894
rect -6454 39658 -6218 39894
rect -6774 39338 -6538 39574
rect -6454 39338 -6218 39574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 8266 708442 8502 708678
rect 8586 708442 8822 708678
rect 8266 708122 8502 708358
rect 8586 708122 8822 708358
rect -5814 669658 -5578 669894
rect -5494 669658 -5258 669894
rect -5814 669338 -5578 669574
rect -5494 669338 -5258 669574
rect -5814 609658 -5578 609894
rect -5494 609658 -5258 609894
rect -5814 609338 -5578 609574
rect -5494 609338 -5258 609574
rect -5814 549658 -5578 549894
rect -5494 549658 -5258 549894
rect -5814 549338 -5578 549574
rect -5494 549338 -5258 549574
rect -5814 489658 -5578 489894
rect -5494 489658 -5258 489894
rect -5814 489338 -5578 489574
rect -5494 489338 -5258 489574
rect -5814 429658 -5578 429894
rect -5494 429658 -5258 429894
rect -5814 429338 -5578 429574
rect -5494 429338 -5258 429574
rect -5814 369658 -5578 369894
rect -5494 369658 -5258 369894
rect -5814 369338 -5578 369574
rect -5494 369338 -5258 369574
rect -5814 309658 -5578 309894
rect -5494 309658 -5258 309894
rect -5814 309338 -5578 309574
rect -5494 309338 -5258 309574
rect -5814 249658 -5578 249894
rect -5494 249658 -5258 249894
rect -5814 249338 -5578 249574
rect -5494 249338 -5258 249574
rect -5814 189658 -5578 189894
rect -5494 189658 -5258 189894
rect -5814 189338 -5578 189574
rect -5494 189338 -5258 189574
rect -5814 129658 -5578 129894
rect -5494 129658 -5258 129894
rect -5814 129338 -5578 129574
rect -5494 129338 -5258 129574
rect -5814 69658 -5578 69894
rect -5494 69658 -5258 69894
rect -5814 69338 -5578 69574
rect -5494 69338 -5258 69574
rect -5814 9658 -5578 9894
rect -5494 9658 -5258 9894
rect -5814 9338 -5578 9574
rect -5494 9338 -5258 9574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 695938 -4618 696174
rect -4534 695938 -4298 696174
rect -4854 695618 -4618 695854
rect -4534 695618 -4298 695854
rect -4854 635938 -4618 636174
rect -4534 635938 -4298 636174
rect -4854 635618 -4618 635854
rect -4534 635618 -4298 635854
rect -4854 575938 -4618 576174
rect -4534 575938 -4298 576174
rect -4854 575618 -4618 575854
rect -4534 575618 -4298 575854
rect -4854 515938 -4618 516174
rect -4534 515938 -4298 516174
rect -4854 515618 -4618 515854
rect -4534 515618 -4298 515854
rect -4854 455938 -4618 456174
rect -4534 455938 -4298 456174
rect -4854 455618 -4618 455854
rect -4534 455618 -4298 455854
rect -4854 395938 -4618 396174
rect -4534 395938 -4298 396174
rect -4854 395618 -4618 395854
rect -4534 395618 -4298 395854
rect -4854 335938 -4618 336174
rect -4534 335938 -4298 336174
rect -4854 335618 -4618 335854
rect -4534 335618 -4298 335854
rect -4854 275938 -4618 276174
rect -4534 275938 -4298 276174
rect -4854 275618 -4618 275854
rect -4534 275618 -4298 275854
rect -4854 215938 -4618 216174
rect -4534 215938 -4298 216174
rect -4854 215618 -4618 215854
rect -4534 215618 -4298 215854
rect -4854 155938 -4618 156174
rect -4534 155938 -4298 156174
rect -4854 155618 -4618 155854
rect -4534 155618 -4298 155854
rect -4854 95938 -4618 96174
rect -4534 95938 -4298 96174
rect -4854 95618 -4618 95854
rect -4534 95618 -4298 95854
rect -4854 35938 -4618 36174
rect -4534 35938 -4298 36174
rect -4854 35618 -4618 35854
rect -4534 35618 -4298 35854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 4546 706522 4782 706758
rect 4866 706522 5102 706758
rect 4546 706202 4782 706438
rect 4866 706202 5102 706438
rect -3894 665938 -3658 666174
rect -3574 665938 -3338 666174
rect -3894 665618 -3658 665854
rect -3574 665618 -3338 665854
rect -3894 605938 -3658 606174
rect -3574 605938 -3338 606174
rect -3894 605618 -3658 605854
rect -3574 605618 -3338 605854
rect -3894 545938 -3658 546174
rect -3574 545938 -3338 546174
rect -3894 545618 -3658 545854
rect -3574 545618 -3338 545854
rect -3894 485938 -3658 486174
rect -3574 485938 -3338 486174
rect -3894 485618 -3658 485854
rect -3574 485618 -3338 485854
rect -3894 425938 -3658 426174
rect -3574 425938 -3338 426174
rect -3894 425618 -3658 425854
rect -3574 425618 -3338 425854
rect -3894 365938 -3658 366174
rect -3574 365938 -3338 366174
rect -3894 365618 -3658 365854
rect -3574 365618 -3338 365854
rect -3894 305938 -3658 306174
rect -3574 305938 -3338 306174
rect -3894 305618 -3658 305854
rect -3574 305618 -3338 305854
rect -3894 245938 -3658 246174
rect -3574 245938 -3338 246174
rect -3894 245618 -3658 245854
rect -3574 245618 -3338 245854
rect -3894 185938 -3658 186174
rect -3574 185938 -3338 186174
rect -3894 185618 -3658 185854
rect -3574 185618 -3338 185854
rect -3894 125938 -3658 126174
rect -3574 125938 -3338 126174
rect -3894 125618 -3658 125854
rect -3574 125618 -3338 125854
rect -3894 65938 -3658 66174
rect -3574 65938 -3338 66174
rect -3894 65618 -3658 65854
rect -3574 65618 -3338 65854
rect -3894 5938 -3658 6174
rect -3574 5938 -3338 6174
rect -3894 5618 -3658 5854
rect -3574 5618 -3338 5854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 692218 -2698 692454
rect -2614 692218 -2378 692454
rect -2934 691898 -2698 692134
rect -2614 691898 -2378 692134
rect -2934 632218 -2698 632454
rect -2614 632218 -2378 632454
rect -2934 631898 -2698 632134
rect -2614 631898 -2378 632134
rect -2934 572218 -2698 572454
rect -2614 572218 -2378 572454
rect -2934 571898 -2698 572134
rect -2614 571898 -2378 572134
rect -2934 512218 -2698 512454
rect -2614 512218 -2378 512454
rect -2934 511898 -2698 512134
rect -2614 511898 -2378 512134
rect -2934 452218 -2698 452454
rect -2614 452218 -2378 452454
rect -2934 451898 -2698 452134
rect -2614 451898 -2378 452134
rect -2934 392218 -2698 392454
rect -2614 392218 -2378 392454
rect -2934 391898 -2698 392134
rect -2614 391898 -2378 392134
rect -2934 332218 -2698 332454
rect -2614 332218 -2378 332454
rect -2934 331898 -2698 332134
rect -2614 331898 -2378 332134
rect -2934 272218 -2698 272454
rect -2614 272218 -2378 272454
rect -2934 271898 -2698 272134
rect -2614 271898 -2378 272134
rect -2934 212218 -2698 212454
rect -2614 212218 -2378 212454
rect -2934 211898 -2698 212134
rect -2614 211898 -2378 212134
rect -2934 152218 -2698 152454
rect -2614 152218 -2378 152454
rect -2934 151898 -2698 152134
rect -2614 151898 -2378 152134
rect -2934 92218 -2698 92454
rect -2614 92218 -2378 92454
rect -2934 91898 -2698 92134
rect -2614 91898 -2378 92134
rect -2934 32218 -2698 32454
rect -2614 32218 -2378 32454
rect -2934 31898 -2698 32134
rect -2614 31898 -2378 32134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 662218 -1738 662454
rect -1654 662218 -1418 662454
rect -1974 661898 -1738 662134
rect -1654 661898 -1418 662134
rect -1974 602218 -1738 602454
rect -1654 602218 -1418 602454
rect -1974 601898 -1738 602134
rect -1654 601898 -1418 602134
rect -1974 542218 -1738 542454
rect -1654 542218 -1418 542454
rect -1974 541898 -1738 542134
rect -1654 541898 -1418 542134
rect -1974 482218 -1738 482454
rect -1654 482218 -1418 482454
rect -1974 481898 -1738 482134
rect -1654 481898 -1418 482134
rect -1974 422218 -1738 422454
rect -1654 422218 -1418 422454
rect -1974 421898 -1738 422134
rect -1654 421898 -1418 422134
rect -1974 362218 -1738 362454
rect -1654 362218 -1418 362454
rect -1974 361898 -1738 362134
rect -1654 361898 -1418 362134
rect -1974 302218 -1738 302454
rect -1654 302218 -1418 302454
rect -1974 301898 -1738 302134
rect -1654 301898 -1418 302134
rect -1974 242218 -1738 242454
rect -1654 242218 -1418 242454
rect -1974 241898 -1738 242134
rect -1654 241898 -1418 242134
rect -1974 182218 -1738 182454
rect -1654 182218 -1418 182454
rect -1974 181898 -1738 182134
rect -1654 181898 -1418 182134
rect -1974 122218 -1738 122454
rect -1654 122218 -1418 122454
rect -1974 121898 -1738 122134
rect -1654 121898 -1418 122134
rect -1974 62218 -1738 62454
rect -1654 62218 -1418 62454
rect -1974 61898 -1738 62134
rect -1654 61898 -1418 62134
rect -1974 2218 -1738 2454
rect -1654 2218 -1418 2454
rect -1974 1898 -1738 2134
rect -1654 1898 -1418 2134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 826 704602 1062 704838
rect 1146 704602 1382 704838
rect 826 704282 1062 704518
rect 1146 704282 1382 704518
rect 826 662218 1062 662454
rect 1146 662218 1382 662454
rect 826 661898 1062 662134
rect 1146 661898 1382 662134
rect 826 602218 1062 602454
rect 1146 602218 1382 602454
rect 826 601898 1062 602134
rect 1146 601898 1382 602134
rect 826 542218 1062 542454
rect 1146 542218 1382 542454
rect 826 541898 1062 542134
rect 1146 541898 1382 542134
rect 826 482218 1062 482454
rect 1146 482218 1382 482454
rect 826 481898 1062 482134
rect 1146 481898 1382 482134
rect 826 422218 1062 422454
rect 1146 422218 1382 422454
rect 826 421898 1062 422134
rect 1146 421898 1382 422134
rect 826 362218 1062 362454
rect 1146 362218 1382 362454
rect 826 361898 1062 362134
rect 1146 361898 1382 362134
rect 4546 665938 4782 666174
rect 4866 665938 5102 666174
rect 4546 665618 4782 665854
rect 4866 665618 5102 665854
rect 4546 605938 4782 606174
rect 4866 605938 5102 606174
rect 4546 605618 4782 605854
rect 4866 605618 5102 605854
rect 4546 545938 4782 546174
rect 4866 545938 5102 546174
rect 4546 545618 4782 545854
rect 4866 545618 5102 545854
rect 4546 485938 4782 486174
rect 4866 485938 5102 486174
rect 4546 485618 4782 485854
rect 4866 485618 5102 485854
rect 4546 425938 4782 426174
rect 4866 425938 5102 426174
rect 4546 425618 4782 425854
rect 4866 425618 5102 425854
rect 4546 365938 4782 366174
rect 4866 365938 5102 366174
rect 4546 365618 4782 365854
rect 4866 365618 5102 365854
rect 826 302218 1062 302454
rect 1146 302218 1382 302454
rect 826 301898 1062 302134
rect 1146 301898 1382 302134
rect 826 242218 1062 242454
rect 1146 242218 1382 242454
rect 826 241898 1062 242134
rect 1146 241898 1382 242134
rect 4546 305938 4782 306174
rect 4866 305938 5102 306174
rect 4546 305618 4782 305854
rect 4866 305618 5102 305854
rect 4546 245938 4782 246174
rect 4866 245938 5102 246174
rect 4546 245618 4782 245854
rect 4866 245618 5102 245854
rect 3286 204222 3522 204458
rect 826 182218 1062 182454
rect 1146 182218 1382 182454
rect 826 181898 1062 182134
rect 1146 181898 1382 182134
rect 826 122218 1062 122454
rect 1146 122218 1382 122454
rect 826 121898 1062 122134
rect 1146 121898 1382 122134
rect 826 62218 1062 62454
rect 1146 62218 1382 62454
rect 826 61898 1062 62134
rect 1146 61898 1382 62134
rect 826 2218 1062 2454
rect 1146 2218 1382 2454
rect 826 1898 1062 2134
rect 1146 1898 1382 2134
rect 826 -582 1062 -346
rect 1146 -582 1382 -346
rect 826 -902 1062 -666
rect 1146 -902 1382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 4546 185938 4782 186174
rect 4866 185938 5102 186174
rect 4546 185618 4782 185854
rect 4866 185618 5102 185854
rect 4546 125938 4782 126174
rect 4866 125938 5102 126174
rect 4546 125618 4782 125854
rect 4866 125618 5102 125854
rect 4546 65938 4782 66174
rect 4866 65938 5102 66174
rect 4546 65618 4782 65854
rect 4866 65618 5102 65854
rect 4546 5938 4782 6174
rect 4866 5938 5102 6174
rect 4546 5618 4782 5854
rect 4866 5618 5102 5854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 4546 -2502 4782 -2266
rect 4866 -2502 5102 -2266
rect 4546 -2822 4782 -2586
rect 4866 -2822 5102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 8266 669658 8502 669894
rect 8586 669658 8822 669894
rect 8266 669338 8502 669574
rect 8586 669338 8822 669574
rect 8266 609658 8502 609894
rect 8586 609658 8822 609894
rect 8266 609338 8502 609574
rect 8586 609338 8822 609574
rect 8266 549658 8502 549894
rect 8586 549658 8822 549894
rect 8266 549338 8502 549574
rect 8586 549338 8822 549574
rect 8266 489658 8502 489894
rect 8586 489658 8822 489894
rect 8266 489338 8502 489574
rect 8586 489338 8822 489574
rect 8266 429658 8502 429894
rect 8586 429658 8822 429894
rect 8266 429338 8502 429574
rect 8586 429338 8822 429574
rect 8266 369658 8502 369894
rect 8586 369658 8822 369894
rect 8266 369338 8502 369574
rect 8586 369338 8822 369574
rect 8266 309658 8502 309894
rect 8586 309658 8822 309894
rect 8266 309338 8502 309574
rect 8586 309338 8822 309574
rect 8266 249658 8502 249894
rect 8586 249658 8822 249894
rect 8266 249338 8502 249574
rect 8586 249338 8822 249574
rect 8266 189658 8502 189894
rect 8586 189658 8822 189894
rect 8266 189338 8502 189574
rect 8586 189338 8822 189574
rect 8266 129658 8502 129894
rect 8586 129658 8822 129894
rect 8266 129338 8502 129574
rect 8586 129338 8822 129574
rect 8266 69658 8502 69894
rect 8586 69658 8822 69894
rect 8266 69338 8502 69574
rect 8586 69338 8822 69574
rect 8266 9658 8502 9894
rect 8586 9658 8822 9894
rect 8266 9338 8502 9574
rect 8586 9338 8822 9574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 8266 -4422 8502 -4186
rect 8586 -4422 8822 -4186
rect 8266 -4742 8502 -4506
rect 8586 -4742 8822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 41986 711322 42222 711558
rect 42306 711322 42542 711558
rect 41986 711002 42222 711238
rect 42306 711002 42542 711238
rect 38266 709402 38502 709638
rect 38586 709402 38822 709638
rect 38266 709082 38502 709318
rect 38586 709082 38822 709318
rect 34546 707482 34782 707718
rect 34866 707482 35102 707718
rect 34546 707162 34782 707398
rect 34866 707162 35102 707398
rect 30826 705562 31062 705798
rect 31146 705562 31382 705798
rect 30826 705242 31062 705478
rect 31146 705242 31382 705478
rect 11986 673378 12222 673614
rect 12306 673378 12542 673614
rect 11986 673058 12222 673294
rect 12306 673058 12542 673294
rect 11986 613378 12222 613614
rect 12306 613378 12542 613614
rect 11986 613058 12222 613294
rect 12306 613058 12542 613294
rect 11986 553378 12222 553614
rect 12306 553378 12542 553614
rect 11986 553058 12222 553294
rect 12306 553058 12542 553294
rect 11986 493378 12222 493614
rect 12306 493378 12542 493614
rect 11986 493058 12222 493294
rect 12306 493058 12542 493294
rect 11986 433378 12222 433614
rect 12306 433378 12542 433614
rect 11986 433058 12222 433294
rect 12306 433058 12542 433294
rect 11986 373378 12222 373614
rect 12306 373378 12542 373614
rect 11986 373058 12222 373294
rect 12306 373058 12542 373294
rect 11986 313378 12222 313614
rect 12306 313378 12542 313614
rect 11986 313058 12222 313294
rect 12306 313058 12542 313294
rect 11986 253378 12222 253614
rect 12306 253378 12542 253614
rect 11986 253058 12222 253294
rect 12306 253058 12542 253294
rect 30826 692218 31062 692454
rect 31146 692218 31382 692454
rect 30826 691898 31062 692134
rect 31146 691898 31382 692134
rect 30826 632218 31062 632454
rect 31146 632218 31382 632454
rect 30826 631898 31062 632134
rect 31146 631898 31382 632134
rect 30826 572218 31062 572454
rect 31146 572218 31382 572454
rect 30826 571898 31062 572134
rect 31146 571898 31382 572134
rect 30826 512218 31062 512454
rect 31146 512218 31382 512454
rect 30826 511898 31062 512134
rect 31146 511898 31382 512134
rect 30826 452218 31062 452454
rect 31146 452218 31382 452454
rect 30826 451898 31062 452134
rect 31146 451898 31382 452134
rect 30826 392218 31062 392454
rect 31146 392218 31382 392454
rect 30826 391898 31062 392134
rect 31146 391898 31382 392134
rect 30826 332218 31062 332454
rect 31146 332218 31382 332454
rect 30826 331898 31062 332134
rect 31146 331898 31382 332134
rect 30826 272218 31062 272454
rect 31146 272218 31382 272454
rect 30826 271898 31062 272134
rect 31146 271898 31382 272134
rect 24630 247062 24866 247298
rect 11986 193378 12222 193614
rect 12306 193378 12542 193614
rect 11986 193058 12222 193294
rect 12306 193058 12542 193294
rect 11986 133378 12222 133614
rect 12306 133378 12542 133614
rect 11986 133058 12222 133294
rect 12306 133058 12542 133294
rect 11986 73378 12222 73614
rect 12306 73378 12542 73614
rect 11986 73058 12222 73294
rect 12306 73058 12542 73294
rect 11986 13378 12222 13614
rect 12306 13378 12542 13614
rect 11986 13058 12222 13294
rect 12306 13058 12542 13294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 30826 212218 31062 212454
rect 31146 212218 31382 212454
rect 30826 211898 31062 212134
rect 31146 211898 31382 212134
rect 30826 152218 31062 152454
rect 31146 152218 31382 152454
rect 30826 151898 31062 152134
rect 31146 151898 31382 152134
rect 30826 92218 31062 92454
rect 31146 92218 31382 92454
rect 30826 91898 31062 92134
rect 31146 91898 31382 92134
rect 30826 32218 31062 32454
rect 31146 32218 31382 32454
rect 30826 31898 31062 32134
rect 31146 31898 31382 32134
rect 30826 -1542 31062 -1306
rect 31146 -1542 31382 -1306
rect 30826 -1862 31062 -1626
rect 31146 -1862 31382 -1626
rect 34546 695938 34782 696174
rect 34866 695938 35102 696174
rect 34546 695618 34782 695854
rect 34866 695618 35102 695854
rect 34546 635938 34782 636174
rect 34866 635938 35102 636174
rect 34546 635618 34782 635854
rect 34866 635618 35102 635854
rect 34546 575938 34782 576174
rect 34866 575938 35102 576174
rect 34546 575618 34782 575854
rect 34866 575618 35102 575854
rect 34546 515938 34782 516174
rect 34866 515938 35102 516174
rect 34546 515618 34782 515854
rect 34866 515618 35102 515854
rect 34546 455938 34782 456174
rect 34866 455938 35102 456174
rect 34546 455618 34782 455854
rect 34866 455618 35102 455854
rect 34546 395938 34782 396174
rect 34866 395938 35102 396174
rect 34546 395618 34782 395854
rect 34866 395618 35102 395854
rect 34546 335938 34782 336174
rect 34866 335938 35102 336174
rect 34546 335618 34782 335854
rect 34866 335618 35102 335854
rect 34546 275938 34782 276174
rect 34866 275938 35102 276174
rect 34546 275618 34782 275854
rect 34866 275618 35102 275854
rect 34546 215938 34782 216174
rect 34866 215938 35102 216174
rect 34546 215618 34782 215854
rect 34866 215618 35102 215854
rect 34546 155938 34782 156174
rect 34866 155938 35102 156174
rect 34546 155618 34782 155854
rect 34866 155618 35102 155854
rect 34546 95938 34782 96174
rect 34866 95938 35102 96174
rect 34546 95618 34782 95854
rect 34866 95618 35102 95854
rect 34546 35938 34782 36174
rect 34866 35938 35102 36174
rect 34546 35618 34782 35854
rect 34866 35618 35102 35854
rect 34546 -3462 34782 -3226
rect 34866 -3462 35102 -3226
rect 34546 -3782 34782 -3546
rect 34866 -3782 35102 -3546
rect 38266 699658 38502 699894
rect 38586 699658 38822 699894
rect 38266 699338 38502 699574
rect 38586 699338 38822 699574
rect 38266 639658 38502 639894
rect 38586 639658 38822 639894
rect 38266 639338 38502 639574
rect 38586 639338 38822 639574
rect 38266 579658 38502 579894
rect 38586 579658 38822 579894
rect 38266 579338 38502 579574
rect 38586 579338 38822 579574
rect 38266 519658 38502 519894
rect 38586 519658 38822 519894
rect 38266 519338 38502 519574
rect 38586 519338 38822 519574
rect 38266 459658 38502 459894
rect 38586 459658 38822 459894
rect 38266 459338 38502 459574
rect 38586 459338 38822 459574
rect 38266 399658 38502 399894
rect 38586 399658 38822 399894
rect 38266 399338 38502 399574
rect 38586 399338 38822 399574
rect 38266 339658 38502 339894
rect 38586 339658 38822 339894
rect 38266 339338 38502 339574
rect 38586 339338 38822 339574
rect 38266 279658 38502 279894
rect 38586 279658 38822 279894
rect 38266 279338 38502 279574
rect 38586 279338 38822 279574
rect 38266 219658 38502 219894
rect 38586 219658 38822 219894
rect 38266 219338 38502 219574
rect 38586 219338 38822 219574
rect 38266 159658 38502 159894
rect 38586 159658 38822 159894
rect 38266 159338 38502 159574
rect 38586 159338 38822 159574
rect 38266 99658 38502 99894
rect 38586 99658 38822 99894
rect 38266 99338 38502 99574
rect 38586 99338 38822 99574
rect 38266 39658 38502 39894
rect 38586 39658 38822 39894
rect 38266 39338 38502 39574
rect 38586 39338 38822 39574
rect 38266 -5382 38502 -5146
rect 38586 -5382 38822 -5146
rect 38266 -5702 38502 -5466
rect 38586 -5702 38822 -5466
rect 71986 710362 72222 710598
rect 72306 710362 72542 710598
rect 71986 710042 72222 710278
rect 72306 710042 72542 710278
rect 68266 708442 68502 708678
rect 68586 708442 68822 708678
rect 68266 708122 68502 708358
rect 68586 708122 68822 708358
rect 64546 706522 64782 706758
rect 64866 706522 65102 706758
rect 64546 706202 64782 706438
rect 64866 706202 65102 706438
rect 41986 643378 42222 643614
rect 42306 643378 42542 643614
rect 41986 643058 42222 643294
rect 42306 643058 42542 643294
rect 41986 583378 42222 583614
rect 42306 583378 42542 583614
rect 41986 583058 42222 583294
rect 42306 583058 42542 583294
rect 41986 523378 42222 523614
rect 42306 523378 42542 523614
rect 41986 523058 42222 523294
rect 42306 523058 42542 523294
rect 41986 463378 42222 463614
rect 42306 463378 42542 463614
rect 41986 463058 42222 463294
rect 42306 463058 42542 463294
rect 41986 403378 42222 403614
rect 42306 403378 42542 403614
rect 41986 403058 42222 403294
rect 42306 403058 42542 403294
rect 41986 343378 42222 343614
rect 42306 343378 42542 343614
rect 41986 343058 42222 343294
rect 42306 343058 42542 343294
rect 41986 283378 42222 283614
rect 42306 283378 42542 283614
rect 41986 283058 42222 283294
rect 42306 283058 42542 283294
rect 41986 223378 42222 223614
rect 42306 223378 42542 223614
rect 41986 223058 42222 223294
rect 42306 223058 42542 223294
rect 41986 163378 42222 163614
rect 42306 163378 42542 163614
rect 41986 163058 42222 163294
rect 42306 163058 42542 163294
rect 41986 103378 42222 103614
rect 42306 103378 42542 103614
rect 41986 103058 42222 103294
rect 42306 103058 42542 103294
rect 41986 43378 42222 43614
rect 42306 43378 42542 43614
rect 41986 43058 42222 43294
rect 42306 43058 42542 43294
rect 11986 -6342 12222 -6106
rect 12306 -6342 12542 -6106
rect 11986 -6662 12222 -6426
rect 12306 -6662 12542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 60826 704602 61062 704838
rect 61146 704602 61382 704838
rect 60826 704282 61062 704518
rect 61146 704282 61382 704518
rect 60826 662218 61062 662454
rect 61146 662218 61382 662454
rect 60826 661898 61062 662134
rect 61146 661898 61382 662134
rect 60826 602218 61062 602454
rect 61146 602218 61382 602454
rect 60826 601898 61062 602134
rect 61146 601898 61382 602134
rect 60826 542218 61062 542454
rect 61146 542218 61382 542454
rect 60826 541898 61062 542134
rect 61146 541898 61382 542134
rect 60826 482218 61062 482454
rect 61146 482218 61382 482454
rect 60826 481898 61062 482134
rect 61146 481898 61382 482134
rect 60826 422218 61062 422454
rect 61146 422218 61382 422454
rect 60826 421898 61062 422134
rect 61146 421898 61382 422134
rect 60826 362218 61062 362454
rect 61146 362218 61382 362454
rect 60826 361898 61062 362134
rect 61146 361898 61382 362134
rect 60826 302218 61062 302454
rect 61146 302218 61382 302454
rect 60826 301898 61062 302134
rect 61146 301898 61382 302134
rect 60826 242218 61062 242454
rect 61146 242218 61382 242454
rect 60826 241898 61062 242134
rect 61146 241898 61382 242134
rect 60826 182218 61062 182454
rect 61146 182218 61382 182454
rect 60826 181898 61062 182134
rect 61146 181898 61382 182134
rect 60826 122218 61062 122454
rect 61146 122218 61382 122454
rect 60826 121898 61062 122134
rect 61146 121898 61382 122134
rect 60826 62218 61062 62454
rect 61146 62218 61382 62454
rect 60826 61898 61062 62134
rect 61146 61898 61382 62134
rect 60826 2218 61062 2454
rect 61146 2218 61382 2454
rect 60826 1898 61062 2134
rect 61146 1898 61382 2134
rect 60826 -582 61062 -346
rect 61146 -582 61382 -346
rect 60826 -902 61062 -666
rect 61146 -902 61382 -666
rect 64546 665938 64782 666174
rect 64866 665938 65102 666174
rect 64546 665618 64782 665854
rect 64866 665618 65102 665854
rect 64546 605938 64782 606174
rect 64866 605938 65102 606174
rect 64546 605618 64782 605854
rect 64866 605618 65102 605854
rect 64546 545938 64782 546174
rect 64866 545938 65102 546174
rect 64546 545618 64782 545854
rect 64866 545618 65102 545854
rect 64546 485938 64782 486174
rect 64866 485938 65102 486174
rect 64546 485618 64782 485854
rect 64866 485618 65102 485854
rect 64546 425938 64782 426174
rect 64866 425938 65102 426174
rect 64546 425618 64782 425854
rect 64866 425618 65102 425854
rect 64546 365938 64782 366174
rect 64866 365938 65102 366174
rect 64546 365618 64782 365854
rect 64866 365618 65102 365854
rect 64546 305938 64782 306174
rect 64866 305938 65102 306174
rect 64546 305618 64782 305854
rect 64866 305618 65102 305854
rect 64546 245938 64782 246174
rect 64866 245938 65102 246174
rect 64546 245618 64782 245854
rect 64866 245618 65102 245854
rect 64546 185938 64782 186174
rect 64866 185938 65102 186174
rect 64546 185618 64782 185854
rect 64866 185618 65102 185854
rect 64546 125938 64782 126174
rect 64866 125938 65102 126174
rect 64546 125618 64782 125854
rect 64866 125618 65102 125854
rect 64546 65938 64782 66174
rect 64866 65938 65102 66174
rect 64546 65618 64782 65854
rect 64866 65618 65102 65854
rect 64546 5938 64782 6174
rect 64866 5938 65102 6174
rect 64546 5618 64782 5854
rect 64866 5618 65102 5854
rect 64546 -2502 64782 -2266
rect 64866 -2502 65102 -2266
rect 64546 -2822 64782 -2586
rect 64866 -2822 65102 -2586
rect 68266 669658 68502 669894
rect 68586 669658 68822 669894
rect 68266 669338 68502 669574
rect 68586 669338 68822 669574
rect 68266 609658 68502 609894
rect 68586 609658 68822 609894
rect 68266 609338 68502 609574
rect 68586 609338 68822 609574
rect 68266 549658 68502 549894
rect 68586 549658 68822 549894
rect 68266 549338 68502 549574
rect 68586 549338 68822 549574
rect 68266 489658 68502 489894
rect 68586 489658 68822 489894
rect 68266 489338 68502 489574
rect 68586 489338 68822 489574
rect 68266 429658 68502 429894
rect 68586 429658 68822 429894
rect 68266 429338 68502 429574
rect 68586 429338 68822 429574
rect 68266 369658 68502 369894
rect 68586 369658 68822 369894
rect 68266 369338 68502 369574
rect 68586 369338 68822 369574
rect 68266 309658 68502 309894
rect 68586 309658 68822 309894
rect 68266 309338 68502 309574
rect 68586 309338 68822 309574
rect 68266 249658 68502 249894
rect 68586 249658 68822 249894
rect 68266 249338 68502 249574
rect 68586 249338 68822 249574
rect 68266 189658 68502 189894
rect 68586 189658 68822 189894
rect 68266 189338 68502 189574
rect 68586 189338 68822 189574
rect 68266 129658 68502 129894
rect 68586 129658 68822 129894
rect 68266 129338 68502 129574
rect 68586 129338 68822 129574
rect 68266 69658 68502 69894
rect 68586 69658 68822 69894
rect 68266 69338 68502 69574
rect 68586 69338 68822 69574
rect 68266 9658 68502 9894
rect 68586 9658 68822 9894
rect 68266 9338 68502 9574
rect 68586 9338 68822 9574
rect 68266 -4422 68502 -4186
rect 68586 -4422 68822 -4186
rect 68266 -4742 68502 -4506
rect 68586 -4742 68822 -4506
rect 101986 711322 102222 711558
rect 102306 711322 102542 711558
rect 101986 711002 102222 711238
rect 102306 711002 102542 711238
rect 98266 709402 98502 709638
rect 98586 709402 98822 709638
rect 98266 709082 98502 709318
rect 98586 709082 98822 709318
rect 94546 707482 94782 707718
rect 94866 707482 95102 707718
rect 94546 707162 94782 707398
rect 94866 707162 95102 707398
rect 71986 673378 72222 673614
rect 72306 673378 72542 673614
rect 71986 673058 72222 673294
rect 72306 673058 72542 673294
rect 71986 613378 72222 613614
rect 72306 613378 72542 613614
rect 71986 613058 72222 613294
rect 72306 613058 72542 613294
rect 71986 553378 72222 553614
rect 72306 553378 72542 553614
rect 71986 553058 72222 553294
rect 72306 553058 72542 553294
rect 71986 493378 72222 493614
rect 72306 493378 72542 493614
rect 71986 493058 72222 493294
rect 72306 493058 72542 493294
rect 71986 433378 72222 433614
rect 72306 433378 72542 433614
rect 71986 433058 72222 433294
rect 72306 433058 72542 433294
rect 71986 373378 72222 373614
rect 72306 373378 72542 373614
rect 71986 373058 72222 373294
rect 72306 373058 72542 373294
rect 71986 313378 72222 313614
rect 72306 313378 72542 313614
rect 71986 313058 72222 313294
rect 72306 313058 72542 313294
rect 71986 253378 72222 253614
rect 72306 253378 72542 253614
rect 71986 253058 72222 253294
rect 72306 253058 72542 253294
rect 71986 193378 72222 193614
rect 72306 193378 72542 193614
rect 71986 193058 72222 193294
rect 72306 193058 72542 193294
rect 71986 133378 72222 133614
rect 72306 133378 72542 133614
rect 71986 133058 72222 133294
rect 72306 133058 72542 133294
rect 71986 73378 72222 73614
rect 72306 73378 72542 73614
rect 71986 73058 72222 73294
rect 72306 73058 72542 73294
rect 71986 13378 72222 13614
rect 72306 13378 72542 13614
rect 71986 13058 72222 13294
rect 72306 13058 72542 13294
rect 41986 -7302 42222 -7066
rect 42306 -7302 42542 -7066
rect 41986 -7622 42222 -7386
rect 42306 -7622 42542 -7386
rect 90826 705562 91062 705798
rect 91146 705562 91382 705798
rect 90826 705242 91062 705478
rect 91146 705242 91382 705478
rect 90826 692218 91062 692454
rect 91146 692218 91382 692454
rect 90826 691898 91062 692134
rect 91146 691898 91382 692134
rect 90826 632218 91062 632454
rect 91146 632218 91382 632454
rect 90826 631898 91062 632134
rect 91146 631898 91382 632134
rect 90826 572218 91062 572454
rect 91146 572218 91382 572454
rect 90826 571898 91062 572134
rect 91146 571898 91382 572134
rect 90826 512218 91062 512454
rect 91146 512218 91382 512454
rect 90826 511898 91062 512134
rect 91146 511898 91382 512134
rect 90826 452218 91062 452454
rect 91146 452218 91382 452454
rect 90826 451898 91062 452134
rect 91146 451898 91382 452134
rect 90826 392218 91062 392454
rect 91146 392218 91382 392454
rect 90826 391898 91062 392134
rect 91146 391898 91382 392134
rect 90826 332218 91062 332454
rect 91146 332218 91382 332454
rect 90826 331898 91062 332134
rect 91146 331898 91382 332134
rect 90826 272218 91062 272454
rect 91146 272218 91382 272454
rect 90826 271898 91062 272134
rect 91146 271898 91382 272134
rect 90826 212218 91062 212454
rect 91146 212218 91382 212454
rect 90826 211898 91062 212134
rect 91146 211898 91382 212134
rect 90826 152218 91062 152454
rect 91146 152218 91382 152454
rect 90826 151898 91062 152134
rect 91146 151898 91382 152134
rect 90826 92218 91062 92454
rect 91146 92218 91382 92454
rect 90826 91898 91062 92134
rect 91146 91898 91382 92134
rect 90826 32218 91062 32454
rect 91146 32218 91382 32454
rect 90826 31898 91062 32134
rect 91146 31898 91382 32134
rect 90826 -1542 91062 -1306
rect 91146 -1542 91382 -1306
rect 90826 -1862 91062 -1626
rect 91146 -1862 91382 -1626
rect 94546 695938 94782 696174
rect 94866 695938 95102 696174
rect 94546 695618 94782 695854
rect 94866 695618 95102 695854
rect 94546 635938 94782 636174
rect 94866 635938 95102 636174
rect 94546 635618 94782 635854
rect 94866 635618 95102 635854
rect 94546 575938 94782 576174
rect 94866 575938 95102 576174
rect 94546 575618 94782 575854
rect 94866 575618 95102 575854
rect 94546 515938 94782 516174
rect 94866 515938 95102 516174
rect 94546 515618 94782 515854
rect 94866 515618 95102 515854
rect 94546 455938 94782 456174
rect 94866 455938 95102 456174
rect 94546 455618 94782 455854
rect 94866 455618 95102 455854
rect 94546 395938 94782 396174
rect 94866 395938 95102 396174
rect 94546 395618 94782 395854
rect 94866 395618 95102 395854
rect 94546 335938 94782 336174
rect 94866 335938 95102 336174
rect 94546 335618 94782 335854
rect 94866 335618 95102 335854
rect 94546 275938 94782 276174
rect 94866 275938 95102 276174
rect 94546 275618 94782 275854
rect 94866 275618 95102 275854
rect 94546 215938 94782 216174
rect 94866 215938 95102 216174
rect 94546 215618 94782 215854
rect 94866 215618 95102 215854
rect 94546 155938 94782 156174
rect 94866 155938 95102 156174
rect 94546 155618 94782 155854
rect 94866 155618 95102 155854
rect 94546 95938 94782 96174
rect 94866 95938 95102 96174
rect 94546 95618 94782 95854
rect 94866 95618 95102 95854
rect 94546 35938 94782 36174
rect 94866 35938 95102 36174
rect 94546 35618 94782 35854
rect 94866 35618 95102 35854
rect 94546 -3462 94782 -3226
rect 94866 -3462 95102 -3226
rect 94546 -3782 94782 -3546
rect 94866 -3782 95102 -3546
rect 98266 699658 98502 699894
rect 98586 699658 98822 699894
rect 98266 699338 98502 699574
rect 98586 699338 98822 699574
rect 98266 639658 98502 639894
rect 98586 639658 98822 639894
rect 98266 639338 98502 639574
rect 98586 639338 98822 639574
rect 98266 579658 98502 579894
rect 98586 579658 98822 579894
rect 98266 579338 98502 579574
rect 98586 579338 98822 579574
rect 98266 519658 98502 519894
rect 98586 519658 98822 519894
rect 98266 519338 98502 519574
rect 98586 519338 98822 519574
rect 98266 459658 98502 459894
rect 98586 459658 98822 459894
rect 98266 459338 98502 459574
rect 98586 459338 98822 459574
rect 98266 399658 98502 399894
rect 98586 399658 98822 399894
rect 98266 399338 98502 399574
rect 98586 399338 98822 399574
rect 98266 339658 98502 339894
rect 98586 339658 98822 339894
rect 98266 339338 98502 339574
rect 98586 339338 98822 339574
rect 98266 279658 98502 279894
rect 98586 279658 98822 279894
rect 98266 279338 98502 279574
rect 98586 279338 98822 279574
rect 98266 219658 98502 219894
rect 98586 219658 98822 219894
rect 98266 219338 98502 219574
rect 98586 219338 98822 219574
rect 98266 159658 98502 159894
rect 98586 159658 98822 159894
rect 98266 159338 98502 159574
rect 98586 159338 98822 159574
rect 98266 99658 98502 99894
rect 98586 99658 98822 99894
rect 98266 99338 98502 99574
rect 98586 99338 98822 99574
rect 98266 39658 98502 39894
rect 98586 39658 98822 39894
rect 98266 39338 98502 39574
rect 98586 39338 98822 39574
rect 98266 -5382 98502 -5146
rect 98586 -5382 98822 -5146
rect 98266 -5702 98502 -5466
rect 98586 -5702 98822 -5466
rect 131986 710362 132222 710598
rect 132306 710362 132542 710598
rect 131986 710042 132222 710278
rect 132306 710042 132542 710278
rect 128266 708442 128502 708678
rect 128586 708442 128822 708678
rect 128266 708122 128502 708358
rect 128586 708122 128822 708358
rect 124546 706522 124782 706758
rect 124866 706522 125102 706758
rect 124546 706202 124782 706438
rect 124866 706202 125102 706438
rect 101986 643378 102222 643614
rect 102306 643378 102542 643614
rect 101986 643058 102222 643294
rect 102306 643058 102542 643294
rect 101986 583378 102222 583614
rect 102306 583378 102542 583614
rect 101986 583058 102222 583294
rect 102306 583058 102542 583294
rect 101986 523378 102222 523614
rect 102306 523378 102542 523614
rect 101986 523058 102222 523294
rect 102306 523058 102542 523294
rect 101986 463378 102222 463614
rect 102306 463378 102542 463614
rect 101986 463058 102222 463294
rect 102306 463058 102542 463294
rect 101986 403378 102222 403614
rect 102306 403378 102542 403614
rect 101986 403058 102222 403294
rect 102306 403058 102542 403294
rect 101986 343378 102222 343614
rect 102306 343378 102542 343614
rect 101986 343058 102222 343294
rect 102306 343058 102542 343294
rect 101986 283378 102222 283614
rect 102306 283378 102542 283614
rect 101986 283058 102222 283294
rect 102306 283058 102542 283294
rect 101986 223378 102222 223614
rect 102306 223378 102542 223614
rect 101986 223058 102222 223294
rect 102306 223058 102542 223294
rect 101986 163378 102222 163614
rect 102306 163378 102542 163614
rect 101986 163058 102222 163294
rect 102306 163058 102542 163294
rect 101986 103378 102222 103614
rect 102306 103378 102542 103614
rect 101986 103058 102222 103294
rect 102306 103058 102542 103294
rect 101986 43378 102222 43614
rect 102306 43378 102542 43614
rect 101986 43058 102222 43294
rect 102306 43058 102542 43294
rect 71986 -6342 72222 -6106
rect 72306 -6342 72542 -6106
rect 71986 -6662 72222 -6426
rect 72306 -6662 72542 -6426
rect 120826 704602 121062 704838
rect 121146 704602 121382 704838
rect 120826 704282 121062 704518
rect 121146 704282 121382 704518
rect 120826 662218 121062 662454
rect 121146 662218 121382 662454
rect 120826 661898 121062 662134
rect 121146 661898 121382 662134
rect 120826 602218 121062 602454
rect 121146 602218 121382 602454
rect 120826 601898 121062 602134
rect 121146 601898 121382 602134
rect 120826 542218 121062 542454
rect 121146 542218 121382 542454
rect 120826 541898 121062 542134
rect 121146 541898 121382 542134
rect 120826 482218 121062 482454
rect 121146 482218 121382 482454
rect 120826 481898 121062 482134
rect 121146 481898 121382 482134
rect 120826 422218 121062 422454
rect 121146 422218 121382 422454
rect 120826 421898 121062 422134
rect 121146 421898 121382 422134
rect 120826 362218 121062 362454
rect 121146 362218 121382 362454
rect 120826 361898 121062 362134
rect 121146 361898 121382 362134
rect 120826 302218 121062 302454
rect 121146 302218 121382 302454
rect 120826 301898 121062 302134
rect 121146 301898 121382 302134
rect 120826 242218 121062 242454
rect 121146 242218 121382 242454
rect 120826 241898 121062 242134
rect 121146 241898 121382 242134
rect 120826 182218 121062 182454
rect 121146 182218 121382 182454
rect 120826 181898 121062 182134
rect 121146 181898 121382 182134
rect 120826 122218 121062 122454
rect 121146 122218 121382 122454
rect 120826 121898 121062 122134
rect 121146 121898 121382 122134
rect 120826 62218 121062 62454
rect 121146 62218 121382 62454
rect 120826 61898 121062 62134
rect 121146 61898 121382 62134
rect 120826 2218 121062 2454
rect 121146 2218 121382 2454
rect 120826 1898 121062 2134
rect 121146 1898 121382 2134
rect 120826 -582 121062 -346
rect 121146 -582 121382 -346
rect 120826 -902 121062 -666
rect 121146 -902 121382 -666
rect 124546 665938 124782 666174
rect 124866 665938 125102 666174
rect 124546 665618 124782 665854
rect 124866 665618 125102 665854
rect 124546 605938 124782 606174
rect 124866 605938 125102 606174
rect 124546 605618 124782 605854
rect 124866 605618 125102 605854
rect 124546 545938 124782 546174
rect 124866 545938 125102 546174
rect 124546 545618 124782 545854
rect 124866 545618 125102 545854
rect 124546 485938 124782 486174
rect 124866 485938 125102 486174
rect 124546 485618 124782 485854
rect 124866 485618 125102 485854
rect 124546 425938 124782 426174
rect 124866 425938 125102 426174
rect 124546 425618 124782 425854
rect 124866 425618 125102 425854
rect 124546 365938 124782 366174
rect 124866 365938 125102 366174
rect 124546 365618 124782 365854
rect 124866 365618 125102 365854
rect 124546 305938 124782 306174
rect 124866 305938 125102 306174
rect 124546 305618 124782 305854
rect 124866 305618 125102 305854
rect 124546 245938 124782 246174
rect 124866 245938 125102 246174
rect 124546 245618 124782 245854
rect 124866 245618 125102 245854
rect 124546 185938 124782 186174
rect 124866 185938 125102 186174
rect 124546 185618 124782 185854
rect 124866 185618 125102 185854
rect 124546 125938 124782 126174
rect 124866 125938 125102 126174
rect 124546 125618 124782 125854
rect 124866 125618 125102 125854
rect 124546 65938 124782 66174
rect 124866 65938 125102 66174
rect 124546 65618 124782 65854
rect 124866 65618 125102 65854
rect 124546 5938 124782 6174
rect 124866 5938 125102 6174
rect 124546 5618 124782 5854
rect 124866 5618 125102 5854
rect 124546 -2502 124782 -2266
rect 124866 -2502 125102 -2266
rect 124546 -2822 124782 -2586
rect 124866 -2822 125102 -2586
rect 128266 669658 128502 669894
rect 128586 669658 128822 669894
rect 128266 669338 128502 669574
rect 128586 669338 128822 669574
rect 128266 609658 128502 609894
rect 128586 609658 128822 609894
rect 128266 609338 128502 609574
rect 128586 609338 128822 609574
rect 128266 549658 128502 549894
rect 128586 549658 128822 549894
rect 128266 549338 128502 549574
rect 128586 549338 128822 549574
rect 128266 489658 128502 489894
rect 128586 489658 128822 489894
rect 128266 489338 128502 489574
rect 128586 489338 128822 489574
rect 128266 429658 128502 429894
rect 128586 429658 128822 429894
rect 128266 429338 128502 429574
rect 128586 429338 128822 429574
rect 128266 369658 128502 369894
rect 128586 369658 128822 369894
rect 128266 369338 128502 369574
rect 128586 369338 128822 369574
rect 128266 309658 128502 309894
rect 128586 309658 128822 309894
rect 128266 309338 128502 309574
rect 128586 309338 128822 309574
rect 128266 249658 128502 249894
rect 128586 249658 128822 249894
rect 128266 249338 128502 249574
rect 128586 249338 128822 249574
rect 128266 189658 128502 189894
rect 128586 189658 128822 189894
rect 128266 189338 128502 189574
rect 128586 189338 128822 189574
rect 128266 129658 128502 129894
rect 128586 129658 128822 129894
rect 128266 129338 128502 129574
rect 128586 129338 128822 129574
rect 128266 69658 128502 69894
rect 128586 69658 128822 69894
rect 128266 69338 128502 69574
rect 128586 69338 128822 69574
rect 128266 9658 128502 9894
rect 128586 9658 128822 9894
rect 128266 9338 128502 9574
rect 128586 9338 128822 9574
rect 128266 -4422 128502 -4186
rect 128586 -4422 128822 -4186
rect 128266 -4742 128502 -4506
rect 128586 -4742 128822 -4506
rect 161986 711322 162222 711558
rect 162306 711322 162542 711558
rect 161986 711002 162222 711238
rect 162306 711002 162542 711238
rect 158266 709402 158502 709638
rect 158586 709402 158822 709638
rect 158266 709082 158502 709318
rect 158586 709082 158822 709318
rect 154546 707482 154782 707718
rect 154866 707482 155102 707718
rect 154546 707162 154782 707398
rect 154866 707162 155102 707398
rect 131986 673378 132222 673614
rect 132306 673378 132542 673614
rect 131986 673058 132222 673294
rect 132306 673058 132542 673294
rect 131986 613378 132222 613614
rect 132306 613378 132542 613614
rect 131986 613058 132222 613294
rect 132306 613058 132542 613294
rect 131986 553378 132222 553614
rect 132306 553378 132542 553614
rect 131986 553058 132222 553294
rect 132306 553058 132542 553294
rect 131986 493378 132222 493614
rect 132306 493378 132542 493614
rect 131986 493058 132222 493294
rect 132306 493058 132542 493294
rect 131986 433378 132222 433614
rect 132306 433378 132542 433614
rect 131986 433058 132222 433294
rect 132306 433058 132542 433294
rect 131986 373378 132222 373614
rect 132306 373378 132542 373614
rect 131986 373058 132222 373294
rect 132306 373058 132542 373294
rect 131986 313378 132222 313614
rect 132306 313378 132542 313614
rect 131986 313058 132222 313294
rect 132306 313058 132542 313294
rect 131986 253378 132222 253614
rect 132306 253378 132542 253614
rect 131986 253058 132222 253294
rect 132306 253058 132542 253294
rect 131986 193378 132222 193614
rect 132306 193378 132542 193614
rect 131986 193058 132222 193294
rect 132306 193058 132542 193294
rect 131986 133378 132222 133614
rect 132306 133378 132542 133614
rect 131986 133058 132222 133294
rect 132306 133058 132542 133294
rect 131986 73378 132222 73614
rect 132306 73378 132542 73614
rect 131986 73058 132222 73294
rect 132306 73058 132542 73294
rect 131986 13378 132222 13614
rect 132306 13378 132542 13614
rect 131986 13058 132222 13294
rect 132306 13058 132542 13294
rect 101986 -7302 102222 -7066
rect 102306 -7302 102542 -7066
rect 101986 -7622 102222 -7386
rect 102306 -7622 102542 -7386
rect 150826 705562 151062 705798
rect 151146 705562 151382 705798
rect 150826 705242 151062 705478
rect 151146 705242 151382 705478
rect 150826 692218 151062 692454
rect 151146 692218 151382 692454
rect 150826 691898 151062 692134
rect 151146 691898 151382 692134
rect 150826 632218 151062 632454
rect 151146 632218 151382 632454
rect 150826 631898 151062 632134
rect 151146 631898 151382 632134
rect 150826 572218 151062 572454
rect 151146 572218 151382 572454
rect 150826 571898 151062 572134
rect 151146 571898 151382 572134
rect 150826 512218 151062 512454
rect 151146 512218 151382 512454
rect 150826 511898 151062 512134
rect 151146 511898 151382 512134
rect 150826 452218 151062 452454
rect 151146 452218 151382 452454
rect 150826 451898 151062 452134
rect 151146 451898 151382 452134
rect 150826 392218 151062 392454
rect 151146 392218 151382 392454
rect 150826 391898 151062 392134
rect 151146 391898 151382 392134
rect 150826 332218 151062 332454
rect 151146 332218 151382 332454
rect 150826 331898 151062 332134
rect 151146 331898 151382 332134
rect 150826 272218 151062 272454
rect 151146 272218 151382 272454
rect 150826 271898 151062 272134
rect 151146 271898 151382 272134
rect 150826 212218 151062 212454
rect 151146 212218 151382 212454
rect 150826 211898 151062 212134
rect 151146 211898 151382 212134
rect 150826 152218 151062 152454
rect 151146 152218 151382 152454
rect 150826 151898 151062 152134
rect 151146 151898 151382 152134
rect 150826 92218 151062 92454
rect 151146 92218 151382 92454
rect 150826 91898 151062 92134
rect 151146 91898 151382 92134
rect 150826 32218 151062 32454
rect 151146 32218 151382 32454
rect 150826 31898 151062 32134
rect 151146 31898 151382 32134
rect 150826 -1542 151062 -1306
rect 151146 -1542 151382 -1306
rect 150826 -1862 151062 -1626
rect 151146 -1862 151382 -1626
rect 154546 695938 154782 696174
rect 154866 695938 155102 696174
rect 154546 695618 154782 695854
rect 154866 695618 155102 695854
rect 154546 635938 154782 636174
rect 154866 635938 155102 636174
rect 154546 635618 154782 635854
rect 154866 635618 155102 635854
rect 154546 575938 154782 576174
rect 154866 575938 155102 576174
rect 154546 575618 154782 575854
rect 154866 575618 155102 575854
rect 154546 515938 154782 516174
rect 154866 515938 155102 516174
rect 154546 515618 154782 515854
rect 154866 515618 155102 515854
rect 154546 455938 154782 456174
rect 154866 455938 155102 456174
rect 154546 455618 154782 455854
rect 154866 455618 155102 455854
rect 154546 395938 154782 396174
rect 154866 395938 155102 396174
rect 154546 395618 154782 395854
rect 154866 395618 155102 395854
rect 154546 335938 154782 336174
rect 154866 335938 155102 336174
rect 154546 335618 154782 335854
rect 154866 335618 155102 335854
rect 154546 275938 154782 276174
rect 154866 275938 155102 276174
rect 154546 275618 154782 275854
rect 154866 275618 155102 275854
rect 154546 215938 154782 216174
rect 154866 215938 155102 216174
rect 154546 215618 154782 215854
rect 154866 215618 155102 215854
rect 154546 155938 154782 156174
rect 154866 155938 155102 156174
rect 154546 155618 154782 155854
rect 154866 155618 155102 155854
rect 154546 95938 154782 96174
rect 154866 95938 155102 96174
rect 154546 95618 154782 95854
rect 154866 95618 155102 95854
rect 154546 35938 154782 36174
rect 154866 35938 155102 36174
rect 154546 35618 154782 35854
rect 154866 35618 155102 35854
rect 154546 -3462 154782 -3226
rect 154866 -3462 155102 -3226
rect 154546 -3782 154782 -3546
rect 154866 -3782 155102 -3546
rect 158266 699658 158502 699894
rect 158586 699658 158822 699894
rect 158266 699338 158502 699574
rect 158586 699338 158822 699574
rect 158266 639658 158502 639894
rect 158586 639658 158822 639894
rect 158266 639338 158502 639574
rect 158586 639338 158822 639574
rect 158266 579658 158502 579894
rect 158586 579658 158822 579894
rect 158266 579338 158502 579574
rect 158586 579338 158822 579574
rect 158266 519658 158502 519894
rect 158586 519658 158822 519894
rect 158266 519338 158502 519574
rect 158586 519338 158822 519574
rect 158266 459658 158502 459894
rect 158586 459658 158822 459894
rect 158266 459338 158502 459574
rect 158586 459338 158822 459574
rect 158266 399658 158502 399894
rect 158586 399658 158822 399894
rect 158266 399338 158502 399574
rect 158586 399338 158822 399574
rect 158266 339658 158502 339894
rect 158586 339658 158822 339894
rect 158266 339338 158502 339574
rect 158586 339338 158822 339574
rect 158266 279658 158502 279894
rect 158586 279658 158822 279894
rect 158266 279338 158502 279574
rect 158586 279338 158822 279574
rect 158266 219658 158502 219894
rect 158586 219658 158822 219894
rect 158266 219338 158502 219574
rect 158586 219338 158822 219574
rect 158266 159658 158502 159894
rect 158586 159658 158822 159894
rect 158266 159338 158502 159574
rect 158586 159338 158822 159574
rect 158266 99658 158502 99894
rect 158586 99658 158822 99894
rect 158266 99338 158502 99574
rect 158586 99338 158822 99574
rect 158266 39658 158502 39894
rect 158586 39658 158822 39894
rect 158266 39338 158502 39574
rect 158586 39338 158822 39574
rect 158266 -5382 158502 -5146
rect 158586 -5382 158822 -5146
rect 158266 -5702 158502 -5466
rect 158586 -5702 158822 -5466
rect 191986 710362 192222 710598
rect 192306 710362 192542 710598
rect 191986 710042 192222 710278
rect 192306 710042 192542 710278
rect 188266 708442 188502 708678
rect 188586 708442 188822 708678
rect 188266 708122 188502 708358
rect 188586 708122 188822 708358
rect 184546 706522 184782 706758
rect 184866 706522 185102 706758
rect 184546 706202 184782 706438
rect 184866 706202 185102 706438
rect 161986 643378 162222 643614
rect 162306 643378 162542 643614
rect 161986 643058 162222 643294
rect 162306 643058 162542 643294
rect 161986 583378 162222 583614
rect 162306 583378 162542 583614
rect 161986 583058 162222 583294
rect 162306 583058 162542 583294
rect 161986 523378 162222 523614
rect 162306 523378 162542 523614
rect 161986 523058 162222 523294
rect 162306 523058 162542 523294
rect 161986 463378 162222 463614
rect 162306 463378 162542 463614
rect 161986 463058 162222 463294
rect 162306 463058 162542 463294
rect 161986 403378 162222 403614
rect 162306 403378 162542 403614
rect 161986 403058 162222 403294
rect 162306 403058 162542 403294
rect 161986 343378 162222 343614
rect 162306 343378 162542 343614
rect 161986 343058 162222 343294
rect 162306 343058 162542 343294
rect 161986 283378 162222 283614
rect 162306 283378 162542 283614
rect 161986 283058 162222 283294
rect 162306 283058 162542 283294
rect 161986 223378 162222 223614
rect 162306 223378 162542 223614
rect 161986 223058 162222 223294
rect 162306 223058 162542 223294
rect 161986 163378 162222 163614
rect 162306 163378 162542 163614
rect 161986 163058 162222 163294
rect 162306 163058 162542 163294
rect 161986 103378 162222 103614
rect 162306 103378 162542 103614
rect 161986 103058 162222 103294
rect 162306 103058 162542 103294
rect 161986 43378 162222 43614
rect 162306 43378 162542 43614
rect 161986 43058 162222 43294
rect 162306 43058 162542 43294
rect 131986 -6342 132222 -6106
rect 132306 -6342 132542 -6106
rect 131986 -6662 132222 -6426
rect 132306 -6662 132542 -6426
rect 180826 704602 181062 704838
rect 181146 704602 181382 704838
rect 180826 704282 181062 704518
rect 181146 704282 181382 704518
rect 180826 662218 181062 662454
rect 181146 662218 181382 662454
rect 180826 661898 181062 662134
rect 181146 661898 181382 662134
rect 180826 602218 181062 602454
rect 181146 602218 181382 602454
rect 180826 601898 181062 602134
rect 181146 601898 181382 602134
rect 180826 542218 181062 542454
rect 181146 542218 181382 542454
rect 180826 541898 181062 542134
rect 181146 541898 181382 542134
rect 180826 482218 181062 482454
rect 181146 482218 181382 482454
rect 180826 481898 181062 482134
rect 181146 481898 181382 482134
rect 180826 422218 181062 422454
rect 181146 422218 181382 422454
rect 180826 421898 181062 422134
rect 181146 421898 181382 422134
rect 180826 362218 181062 362454
rect 181146 362218 181382 362454
rect 180826 361898 181062 362134
rect 181146 361898 181382 362134
rect 180826 302218 181062 302454
rect 181146 302218 181382 302454
rect 180826 301898 181062 302134
rect 181146 301898 181382 302134
rect 180826 242218 181062 242454
rect 181146 242218 181382 242454
rect 180826 241898 181062 242134
rect 181146 241898 181382 242134
rect 180826 182218 181062 182454
rect 181146 182218 181382 182454
rect 180826 181898 181062 182134
rect 181146 181898 181382 182134
rect 180826 122218 181062 122454
rect 181146 122218 181382 122454
rect 180826 121898 181062 122134
rect 181146 121898 181382 122134
rect 180826 62218 181062 62454
rect 181146 62218 181382 62454
rect 180826 61898 181062 62134
rect 181146 61898 181382 62134
rect 180826 2218 181062 2454
rect 181146 2218 181382 2454
rect 180826 1898 181062 2134
rect 181146 1898 181382 2134
rect 180826 -582 181062 -346
rect 181146 -582 181382 -346
rect 180826 -902 181062 -666
rect 181146 -902 181382 -666
rect 184546 665938 184782 666174
rect 184866 665938 185102 666174
rect 184546 665618 184782 665854
rect 184866 665618 185102 665854
rect 184546 605938 184782 606174
rect 184866 605938 185102 606174
rect 184546 605618 184782 605854
rect 184866 605618 185102 605854
rect 184546 545938 184782 546174
rect 184866 545938 185102 546174
rect 184546 545618 184782 545854
rect 184866 545618 185102 545854
rect 184546 485938 184782 486174
rect 184866 485938 185102 486174
rect 184546 485618 184782 485854
rect 184866 485618 185102 485854
rect 184546 425938 184782 426174
rect 184866 425938 185102 426174
rect 184546 425618 184782 425854
rect 184866 425618 185102 425854
rect 184546 365938 184782 366174
rect 184866 365938 185102 366174
rect 184546 365618 184782 365854
rect 184866 365618 185102 365854
rect 184546 305938 184782 306174
rect 184866 305938 185102 306174
rect 184546 305618 184782 305854
rect 184866 305618 185102 305854
rect 184546 245938 184782 246174
rect 184866 245938 185102 246174
rect 184546 245618 184782 245854
rect 184866 245618 185102 245854
rect 184546 185938 184782 186174
rect 184866 185938 185102 186174
rect 184546 185618 184782 185854
rect 184866 185618 185102 185854
rect 184546 125938 184782 126174
rect 184866 125938 185102 126174
rect 184546 125618 184782 125854
rect 184866 125618 185102 125854
rect 184546 65938 184782 66174
rect 184866 65938 185102 66174
rect 184546 65618 184782 65854
rect 184866 65618 185102 65854
rect 184546 5938 184782 6174
rect 184866 5938 185102 6174
rect 184546 5618 184782 5854
rect 184866 5618 185102 5854
rect 184546 -2502 184782 -2266
rect 184866 -2502 185102 -2266
rect 184546 -2822 184782 -2586
rect 184866 -2822 185102 -2586
rect 188266 669658 188502 669894
rect 188586 669658 188822 669894
rect 188266 669338 188502 669574
rect 188586 669338 188822 669574
rect 188266 609658 188502 609894
rect 188586 609658 188822 609894
rect 188266 609338 188502 609574
rect 188586 609338 188822 609574
rect 188266 549658 188502 549894
rect 188586 549658 188822 549894
rect 188266 549338 188502 549574
rect 188586 549338 188822 549574
rect 188266 489658 188502 489894
rect 188586 489658 188822 489894
rect 188266 489338 188502 489574
rect 188586 489338 188822 489574
rect 188266 429658 188502 429894
rect 188586 429658 188822 429894
rect 188266 429338 188502 429574
rect 188586 429338 188822 429574
rect 188266 369658 188502 369894
rect 188586 369658 188822 369894
rect 188266 369338 188502 369574
rect 188586 369338 188822 369574
rect 188266 309658 188502 309894
rect 188586 309658 188822 309894
rect 188266 309338 188502 309574
rect 188586 309338 188822 309574
rect 188266 249658 188502 249894
rect 188586 249658 188822 249894
rect 188266 249338 188502 249574
rect 188586 249338 188822 249574
rect 188266 189658 188502 189894
rect 188586 189658 188822 189894
rect 188266 189338 188502 189574
rect 188586 189338 188822 189574
rect 188266 129658 188502 129894
rect 188586 129658 188822 129894
rect 188266 129338 188502 129574
rect 188586 129338 188822 129574
rect 188266 69658 188502 69894
rect 188586 69658 188822 69894
rect 188266 69338 188502 69574
rect 188586 69338 188822 69574
rect 188266 9658 188502 9894
rect 188586 9658 188822 9894
rect 188266 9338 188502 9574
rect 188586 9338 188822 9574
rect 188266 -4422 188502 -4186
rect 188586 -4422 188822 -4186
rect 188266 -4742 188502 -4506
rect 188586 -4742 188822 -4506
rect 221986 711322 222222 711558
rect 222306 711322 222542 711558
rect 221986 711002 222222 711238
rect 222306 711002 222542 711238
rect 218266 709402 218502 709638
rect 218586 709402 218822 709638
rect 218266 709082 218502 709318
rect 218586 709082 218822 709318
rect 214546 707482 214782 707718
rect 214866 707482 215102 707718
rect 214546 707162 214782 707398
rect 214866 707162 215102 707398
rect 191986 673378 192222 673614
rect 192306 673378 192542 673614
rect 191986 673058 192222 673294
rect 192306 673058 192542 673294
rect 191986 613378 192222 613614
rect 192306 613378 192542 613614
rect 191986 613058 192222 613294
rect 192306 613058 192542 613294
rect 191986 553378 192222 553614
rect 192306 553378 192542 553614
rect 191986 553058 192222 553294
rect 192306 553058 192542 553294
rect 191986 493378 192222 493614
rect 192306 493378 192542 493614
rect 191986 493058 192222 493294
rect 192306 493058 192542 493294
rect 191986 433378 192222 433614
rect 192306 433378 192542 433614
rect 191986 433058 192222 433294
rect 192306 433058 192542 433294
rect 191986 373378 192222 373614
rect 192306 373378 192542 373614
rect 191986 373058 192222 373294
rect 192306 373058 192542 373294
rect 191986 313378 192222 313614
rect 192306 313378 192542 313614
rect 191986 313058 192222 313294
rect 192306 313058 192542 313294
rect 210826 705562 211062 705798
rect 211146 705562 211382 705798
rect 210826 705242 211062 705478
rect 211146 705242 211382 705478
rect 210826 692218 211062 692454
rect 211146 692218 211382 692454
rect 210826 691898 211062 692134
rect 211146 691898 211382 692134
rect 210826 632218 211062 632454
rect 211146 632218 211382 632454
rect 210826 631898 211062 632134
rect 211146 631898 211382 632134
rect 210826 572218 211062 572454
rect 211146 572218 211382 572454
rect 210826 571898 211062 572134
rect 211146 571898 211382 572134
rect 210826 512218 211062 512454
rect 211146 512218 211382 512454
rect 210826 511898 211062 512134
rect 211146 511898 211382 512134
rect 210826 452218 211062 452454
rect 211146 452218 211382 452454
rect 210826 451898 211062 452134
rect 211146 451898 211382 452134
rect 210826 392218 211062 392454
rect 211146 392218 211382 392454
rect 210826 391898 211062 392134
rect 211146 391898 211382 392134
rect 210826 332218 211062 332454
rect 211146 332218 211382 332454
rect 210826 331898 211062 332134
rect 211146 331898 211382 332134
rect 210826 272218 211062 272454
rect 211146 272218 211382 272454
rect 210826 271898 211062 272134
rect 211146 271898 211382 272134
rect 214546 695938 214782 696174
rect 214866 695938 215102 696174
rect 214546 695618 214782 695854
rect 214866 695618 215102 695854
rect 214546 635938 214782 636174
rect 214866 635938 215102 636174
rect 214546 635618 214782 635854
rect 214866 635618 215102 635854
rect 214546 575938 214782 576174
rect 214866 575938 215102 576174
rect 214546 575618 214782 575854
rect 214866 575618 215102 575854
rect 214546 515938 214782 516174
rect 214866 515938 215102 516174
rect 214546 515618 214782 515854
rect 214866 515618 215102 515854
rect 214546 455938 214782 456174
rect 214866 455938 215102 456174
rect 214546 455618 214782 455854
rect 214866 455618 215102 455854
rect 214546 395938 214782 396174
rect 214866 395938 215102 396174
rect 214546 395618 214782 395854
rect 214866 395618 215102 395854
rect 214546 335938 214782 336174
rect 214866 335938 215102 336174
rect 214546 335618 214782 335854
rect 214866 335618 215102 335854
rect 214546 275938 214782 276174
rect 214866 275938 215102 276174
rect 214546 275618 214782 275854
rect 214866 275618 215102 275854
rect 218266 699658 218502 699894
rect 218586 699658 218822 699894
rect 218266 699338 218502 699574
rect 218586 699338 218822 699574
rect 218266 639658 218502 639894
rect 218586 639658 218822 639894
rect 218266 639338 218502 639574
rect 218586 639338 218822 639574
rect 218266 579658 218502 579894
rect 218586 579658 218822 579894
rect 218266 579338 218502 579574
rect 218586 579338 218822 579574
rect 218266 519658 218502 519894
rect 218586 519658 218822 519894
rect 218266 519338 218502 519574
rect 218586 519338 218822 519574
rect 218266 459658 218502 459894
rect 218586 459658 218822 459894
rect 218266 459338 218502 459574
rect 218586 459338 218822 459574
rect 218266 399658 218502 399894
rect 218586 399658 218822 399894
rect 218266 399338 218502 399574
rect 218586 399338 218822 399574
rect 218266 339658 218502 339894
rect 218586 339658 218822 339894
rect 218266 339338 218502 339574
rect 218586 339338 218822 339574
rect 218266 279658 218502 279894
rect 218586 279658 218822 279894
rect 218266 279338 218502 279574
rect 218586 279338 218822 279574
rect 191986 253378 192222 253614
rect 192306 253378 192542 253614
rect 191986 253058 192222 253294
rect 192306 253058 192542 253294
rect 204250 242218 204486 242454
rect 204250 241898 204486 242134
rect 191986 193378 192222 193614
rect 192306 193378 192542 193614
rect 191986 193058 192222 193294
rect 192306 193058 192542 193294
rect 191986 133378 192222 133614
rect 192306 133378 192542 133614
rect 191986 133058 192222 133294
rect 192306 133058 192542 133294
rect 191986 73378 192222 73614
rect 192306 73378 192542 73614
rect 191986 73058 192222 73294
rect 192306 73058 192542 73294
rect 191986 13378 192222 13614
rect 192306 13378 192542 13614
rect 191986 13058 192222 13294
rect 192306 13058 192542 13294
rect 161986 -7302 162222 -7066
rect 162306 -7302 162542 -7066
rect 161986 -7622 162222 -7386
rect 162306 -7622 162542 -7386
rect 251986 710362 252222 710598
rect 252306 710362 252542 710598
rect 251986 710042 252222 710278
rect 252306 710042 252542 710278
rect 248266 708442 248502 708678
rect 248586 708442 248822 708678
rect 248266 708122 248502 708358
rect 248586 708122 248822 708358
rect 244546 706522 244782 706758
rect 244866 706522 245102 706758
rect 244546 706202 244782 706438
rect 244866 706202 245102 706438
rect 221986 643378 222222 643614
rect 222306 643378 222542 643614
rect 221986 643058 222222 643294
rect 222306 643058 222542 643294
rect 221986 583378 222222 583614
rect 222306 583378 222542 583614
rect 221986 583058 222222 583294
rect 222306 583058 222542 583294
rect 221986 523378 222222 523614
rect 222306 523378 222542 523614
rect 221986 523058 222222 523294
rect 222306 523058 222542 523294
rect 221986 463378 222222 463614
rect 222306 463378 222542 463614
rect 221986 463058 222222 463294
rect 222306 463058 222542 463294
rect 221986 403378 222222 403614
rect 222306 403378 222542 403614
rect 221986 403058 222222 403294
rect 222306 403058 222542 403294
rect 221986 343378 222222 343614
rect 222306 343378 222542 343614
rect 221986 343058 222222 343294
rect 222306 343058 222542 343294
rect 221986 283378 222222 283614
rect 222306 283378 222542 283614
rect 221986 283058 222222 283294
rect 222306 283058 222542 283294
rect 240826 704602 241062 704838
rect 241146 704602 241382 704838
rect 240826 704282 241062 704518
rect 241146 704282 241382 704518
rect 240826 662218 241062 662454
rect 241146 662218 241382 662454
rect 240826 661898 241062 662134
rect 241146 661898 241382 662134
rect 240826 602218 241062 602454
rect 241146 602218 241382 602454
rect 240826 601898 241062 602134
rect 241146 601898 241382 602134
rect 240826 542218 241062 542454
rect 241146 542218 241382 542454
rect 240826 541898 241062 542134
rect 241146 541898 241382 542134
rect 240826 482218 241062 482454
rect 241146 482218 241382 482454
rect 240826 481898 241062 482134
rect 241146 481898 241382 482134
rect 240826 422218 241062 422454
rect 241146 422218 241382 422454
rect 240826 421898 241062 422134
rect 241146 421898 241382 422134
rect 240826 362218 241062 362454
rect 241146 362218 241382 362454
rect 240826 361898 241062 362134
rect 241146 361898 241382 362134
rect 240826 302218 241062 302454
rect 241146 302218 241382 302454
rect 240826 301898 241062 302134
rect 241146 301898 241382 302134
rect 244546 665938 244782 666174
rect 244866 665938 245102 666174
rect 244546 665618 244782 665854
rect 244866 665618 245102 665854
rect 244546 605938 244782 606174
rect 244866 605938 245102 606174
rect 244546 605618 244782 605854
rect 244866 605618 245102 605854
rect 244546 545938 244782 546174
rect 244866 545938 245102 546174
rect 244546 545618 244782 545854
rect 244866 545618 245102 545854
rect 244546 485938 244782 486174
rect 244866 485938 245102 486174
rect 244546 485618 244782 485854
rect 244866 485618 245102 485854
rect 244546 425938 244782 426174
rect 244866 425938 245102 426174
rect 244546 425618 244782 425854
rect 244866 425618 245102 425854
rect 244546 365938 244782 366174
rect 244866 365938 245102 366174
rect 244546 365618 244782 365854
rect 244866 365618 245102 365854
rect 244546 305938 244782 306174
rect 244866 305938 245102 306174
rect 244546 305618 244782 305854
rect 244866 305618 245102 305854
rect 248266 669658 248502 669894
rect 248586 669658 248822 669894
rect 248266 669338 248502 669574
rect 248586 669338 248822 669574
rect 248266 609658 248502 609894
rect 248586 609658 248822 609894
rect 248266 609338 248502 609574
rect 248586 609338 248822 609574
rect 248266 549658 248502 549894
rect 248586 549658 248822 549894
rect 248266 549338 248502 549574
rect 248586 549338 248822 549574
rect 248266 489658 248502 489894
rect 248586 489658 248822 489894
rect 248266 489338 248502 489574
rect 248586 489338 248822 489574
rect 248266 429658 248502 429894
rect 248586 429658 248822 429894
rect 248266 429338 248502 429574
rect 248586 429338 248822 429574
rect 248266 369658 248502 369894
rect 248586 369658 248822 369894
rect 248266 369338 248502 369574
rect 248586 369338 248822 369574
rect 248266 309658 248502 309894
rect 248586 309658 248822 309894
rect 248266 309338 248502 309574
rect 248586 309338 248822 309574
rect 281986 711322 282222 711558
rect 282306 711322 282542 711558
rect 281986 711002 282222 711238
rect 282306 711002 282542 711238
rect 278266 709402 278502 709638
rect 278586 709402 278822 709638
rect 278266 709082 278502 709318
rect 278586 709082 278822 709318
rect 274546 707482 274782 707718
rect 274866 707482 275102 707718
rect 274546 707162 274782 707398
rect 274866 707162 275102 707398
rect 251986 673378 252222 673614
rect 252306 673378 252542 673614
rect 251986 673058 252222 673294
rect 252306 673058 252542 673294
rect 251986 613378 252222 613614
rect 252306 613378 252542 613614
rect 251986 613058 252222 613294
rect 252306 613058 252542 613294
rect 251986 553378 252222 553614
rect 252306 553378 252542 553614
rect 251986 553058 252222 553294
rect 252306 553058 252542 553294
rect 251986 493378 252222 493614
rect 252306 493378 252542 493614
rect 251986 493058 252222 493294
rect 252306 493058 252542 493294
rect 251986 433378 252222 433614
rect 252306 433378 252542 433614
rect 251986 433058 252222 433294
rect 252306 433058 252542 433294
rect 251986 373378 252222 373614
rect 252306 373378 252542 373614
rect 251986 373058 252222 373294
rect 252306 373058 252542 373294
rect 251986 313378 252222 313614
rect 252306 313378 252542 313614
rect 251986 313058 252222 313294
rect 252306 313058 252542 313294
rect 270826 705562 271062 705798
rect 271146 705562 271382 705798
rect 270826 705242 271062 705478
rect 271146 705242 271382 705478
rect 270826 692218 271062 692454
rect 271146 692218 271382 692454
rect 270826 691898 271062 692134
rect 271146 691898 271382 692134
rect 270826 632218 271062 632454
rect 271146 632218 271382 632454
rect 270826 631898 271062 632134
rect 271146 631898 271382 632134
rect 270826 572218 271062 572454
rect 271146 572218 271382 572454
rect 270826 571898 271062 572134
rect 271146 571898 271382 572134
rect 270826 512218 271062 512454
rect 271146 512218 271382 512454
rect 270826 511898 271062 512134
rect 271146 511898 271382 512134
rect 270826 452218 271062 452454
rect 271146 452218 271382 452454
rect 270826 451898 271062 452134
rect 271146 451898 271382 452134
rect 270826 392218 271062 392454
rect 271146 392218 271382 392454
rect 270826 391898 271062 392134
rect 271146 391898 271382 392134
rect 270826 332218 271062 332454
rect 271146 332218 271382 332454
rect 270826 331898 271062 332134
rect 271146 331898 271382 332134
rect 270826 272218 271062 272454
rect 271146 272218 271382 272454
rect 270826 271898 271062 272134
rect 271146 271898 271382 272134
rect 249478 247062 249714 247298
rect 234970 242218 235206 242454
rect 234970 241898 235206 242134
rect 218198 217822 218434 218058
rect 249478 217822 249714 218058
rect 219610 212218 219846 212454
rect 219610 211898 219846 212134
rect 270826 212218 271062 212454
rect 271146 212218 271382 212454
rect 270826 211898 271062 212134
rect 271146 211898 271382 212134
rect 249478 204222 249714 204458
rect 210826 152218 211062 152454
rect 211146 152218 211382 152454
rect 210826 151898 211062 152134
rect 211146 151898 211382 152134
rect 210826 92218 211062 92454
rect 211146 92218 211382 92454
rect 210826 91898 211062 92134
rect 211146 91898 211382 92134
rect 210826 32218 211062 32454
rect 211146 32218 211382 32454
rect 210826 31898 211062 32134
rect 211146 31898 211382 32134
rect 210826 -1542 211062 -1306
rect 211146 -1542 211382 -1306
rect 210826 -1862 211062 -1626
rect 211146 -1862 211382 -1626
rect 214546 155938 214782 156174
rect 214866 155938 215102 156174
rect 214546 155618 214782 155854
rect 214866 155618 215102 155854
rect 214546 95938 214782 96174
rect 214866 95938 215102 96174
rect 214546 95618 214782 95854
rect 214866 95618 215102 95854
rect 214546 35938 214782 36174
rect 214866 35938 215102 36174
rect 214546 35618 214782 35854
rect 214866 35618 215102 35854
rect 214546 -3462 214782 -3226
rect 214866 -3462 215102 -3226
rect 214546 -3782 214782 -3546
rect 214866 -3782 215102 -3546
rect 218266 159658 218502 159894
rect 218586 159658 218822 159894
rect 218266 159338 218502 159574
rect 218586 159338 218822 159574
rect 218266 99658 218502 99894
rect 218586 99658 218822 99894
rect 218266 99338 218502 99574
rect 218586 99338 218822 99574
rect 218266 39658 218502 39894
rect 218586 39658 218822 39894
rect 218266 39338 218502 39574
rect 218586 39338 218822 39574
rect 218266 -5382 218502 -5146
rect 218586 -5382 218822 -5146
rect 218266 -5702 218502 -5466
rect 218586 -5702 218822 -5466
rect 221986 163378 222222 163614
rect 222306 163378 222542 163614
rect 221986 163058 222222 163294
rect 222306 163058 222542 163294
rect 221986 103378 222222 103614
rect 222306 103378 222542 103614
rect 221986 103058 222222 103294
rect 222306 103058 222542 103294
rect 221986 43378 222222 43614
rect 222306 43378 222542 43614
rect 221986 43058 222222 43294
rect 222306 43058 222542 43294
rect 191986 -6342 192222 -6106
rect 192306 -6342 192542 -6106
rect 191986 -6662 192222 -6426
rect 192306 -6662 192542 -6426
rect 240826 182218 241062 182454
rect 241146 182218 241382 182454
rect 240826 181898 241062 182134
rect 241146 181898 241382 182134
rect 240826 122218 241062 122454
rect 241146 122218 241382 122454
rect 240826 121898 241062 122134
rect 241146 121898 241382 122134
rect 240826 62218 241062 62454
rect 241146 62218 241382 62454
rect 240826 61898 241062 62134
rect 241146 61898 241382 62134
rect 240826 2218 241062 2454
rect 241146 2218 241382 2454
rect 240826 1898 241062 2134
rect 241146 1898 241382 2134
rect 240826 -582 241062 -346
rect 241146 -582 241382 -346
rect 240826 -902 241062 -666
rect 241146 -902 241382 -666
rect 244546 185938 244782 186174
rect 244866 185938 245102 186174
rect 244546 185618 244782 185854
rect 244866 185618 245102 185854
rect 244546 125938 244782 126174
rect 244866 125938 245102 126174
rect 244546 125618 244782 125854
rect 244866 125618 245102 125854
rect 244546 65938 244782 66174
rect 244866 65938 245102 66174
rect 244546 65618 244782 65854
rect 244866 65618 245102 65854
rect 244546 5938 244782 6174
rect 244866 5938 245102 6174
rect 244546 5618 244782 5854
rect 244866 5618 245102 5854
rect 244546 -2502 244782 -2266
rect 244866 -2502 245102 -2266
rect 244546 -2822 244782 -2586
rect 244866 -2822 245102 -2586
rect 248266 189658 248502 189894
rect 248586 189658 248822 189894
rect 248266 189338 248502 189574
rect 248586 189338 248822 189574
rect 248266 129658 248502 129894
rect 248586 129658 248822 129894
rect 248266 129338 248502 129574
rect 248586 129338 248822 129574
rect 248266 69658 248502 69894
rect 248586 69658 248822 69894
rect 248266 69338 248502 69574
rect 248586 69338 248822 69574
rect 248266 9658 248502 9894
rect 248586 9658 248822 9894
rect 248266 9338 248502 9574
rect 248586 9338 248822 9574
rect 248266 -4422 248502 -4186
rect 248586 -4422 248822 -4186
rect 248266 -4742 248502 -4506
rect 248586 -4742 248822 -4506
rect 251986 193378 252222 193614
rect 252306 193378 252542 193614
rect 251986 193058 252222 193294
rect 252306 193058 252542 193294
rect 251986 133378 252222 133614
rect 252306 133378 252542 133614
rect 251986 133058 252222 133294
rect 252306 133058 252542 133294
rect 251986 73378 252222 73614
rect 252306 73378 252542 73614
rect 251986 73058 252222 73294
rect 252306 73058 252542 73294
rect 251986 13378 252222 13614
rect 252306 13378 252542 13614
rect 251986 13058 252222 13294
rect 252306 13058 252542 13294
rect 221986 -7302 222222 -7066
rect 222306 -7302 222542 -7066
rect 221986 -7622 222222 -7386
rect 222306 -7622 222542 -7386
rect 270826 152218 271062 152454
rect 271146 152218 271382 152454
rect 270826 151898 271062 152134
rect 271146 151898 271382 152134
rect 270826 92218 271062 92454
rect 271146 92218 271382 92454
rect 270826 91898 271062 92134
rect 271146 91898 271382 92134
rect 270826 32218 271062 32454
rect 271146 32218 271382 32454
rect 270826 31898 271062 32134
rect 271146 31898 271382 32134
rect 270826 -1542 271062 -1306
rect 271146 -1542 271382 -1306
rect 270826 -1862 271062 -1626
rect 271146 -1862 271382 -1626
rect 274546 695938 274782 696174
rect 274866 695938 275102 696174
rect 274546 695618 274782 695854
rect 274866 695618 275102 695854
rect 274546 635938 274782 636174
rect 274866 635938 275102 636174
rect 274546 635618 274782 635854
rect 274866 635618 275102 635854
rect 274546 575938 274782 576174
rect 274866 575938 275102 576174
rect 274546 575618 274782 575854
rect 274866 575618 275102 575854
rect 274546 515938 274782 516174
rect 274866 515938 275102 516174
rect 274546 515618 274782 515854
rect 274866 515618 275102 515854
rect 274546 455938 274782 456174
rect 274866 455938 275102 456174
rect 274546 455618 274782 455854
rect 274866 455618 275102 455854
rect 274546 395938 274782 396174
rect 274866 395938 275102 396174
rect 274546 395618 274782 395854
rect 274866 395618 275102 395854
rect 274546 335938 274782 336174
rect 274866 335938 275102 336174
rect 274546 335618 274782 335854
rect 274866 335618 275102 335854
rect 274546 275938 274782 276174
rect 274866 275938 275102 276174
rect 274546 275618 274782 275854
rect 274866 275618 275102 275854
rect 274546 215938 274782 216174
rect 274866 215938 275102 216174
rect 274546 215618 274782 215854
rect 274866 215618 275102 215854
rect 274546 155938 274782 156174
rect 274866 155938 275102 156174
rect 274546 155618 274782 155854
rect 274866 155618 275102 155854
rect 274546 95938 274782 96174
rect 274866 95938 275102 96174
rect 274546 95618 274782 95854
rect 274866 95618 275102 95854
rect 274546 35938 274782 36174
rect 274866 35938 275102 36174
rect 274546 35618 274782 35854
rect 274866 35618 275102 35854
rect 274546 -3462 274782 -3226
rect 274866 -3462 275102 -3226
rect 274546 -3782 274782 -3546
rect 274866 -3782 275102 -3546
rect 278266 699658 278502 699894
rect 278586 699658 278822 699894
rect 278266 699338 278502 699574
rect 278586 699338 278822 699574
rect 278266 639658 278502 639894
rect 278586 639658 278822 639894
rect 278266 639338 278502 639574
rect 278586 639338 278822 639574
rect 278266 579658 278502 579894
rect 278586 579658 278822 579894
rect 278266 579338 278502 579574
rect 278586 579338 278822 579574
rect 278266 519658 278502 519894
rect 278586 519658 278822 519894
rect 278266 519338 278502 519574
rect 278586 519338 278822 519574
rect 278266 459658 278502 459894
rect 278586 459658 278822 459894
rect 278266 459338 278502 459574
rect 278586 459338 278822 459574
rect 278266 399658 278502 399894
rect 278586 399658 278822 399894
rect 278266 399338 278502 399574
rect 278586 399338 278822 399574
rect 278266 339658 278502 339894
rect 278586 339658 278822 339894
rect 278266 339338 278502 339574
rect 278586 339338 278822 339574
rect 278266 279658 278502 279894
rect 278586 279658 278822 279894
rect 278266 279338 278502 279574
rect 278586 279338 278822 279574
rect 278266 219658 278502 219894
rect 278586 219658 278822 219894
rect 278266 219338 278502 219574
rect 278586 219338 278822 219574
rect 278266 159658 278502 159894
rect 278586 159658 278822 159894
rect 278266 159338 278502 159574
rect 278586 159338 278822 159574
rect 278266 99658 278502 99894
rect 278586 99658 278822 99894
rect 278266 99338 278502 99574
rect 278586 99338 278822 99574
rect 278266 39658 278502 39894
rect 278586 39658 278822 39894
rect 278266 39338 278502 39574
rect 278586 39338 278822 39574
rect 278266 -5382 278502 -5146
rect 278586 -5382 278822 -5146
rect 278266 -5702 278502 -5466
rect 278586 -5702 278822 -5466
rect 311986 710362 312222 710598
rect 312306 710362 312542 710598
rect 311986 710042 312222 710278
rect 312306 710042 312542 710278
rect 308266 708442 308502 708678
rect 308586 708442 308822 708678
rect 308266 708122 308502 708358
rect 308586 708122 308822 708358
rect 304546 706522 304782 706758
rect 304866 706522 305102 706758
rect 304546 706202 304782 706438
rect 304866 706202 305102 706438
rect 281986 643378 282222 643614
rect 282306 643378 282542 643614
rect 281986 643058 282222 643294
rect 282306 643058 282542 643294
rect 281986 583378 282222 583614
rect 282306 583378 282542 583614
rect 281986 583058 282222 583294
rect 282306 583058 282542 583294
rect 281986 523378 282222 523614
rect 282306 523378 282542 523614
rect 281986 523058 282222 523294
rect 282306 523058 282542 523294
rect 281986 463378 282222 463614
rect 282306 463378 282542 463614
rect 281986 463058 282222 463294
rect 282306 463058 282542 463294
rect 281986 403378 282222 403614
rect 282306 403378 282542 403614
rect 281986 403058 282222 403294
rect 282306 403058 282542 403294
rect 281986 343378 282222 343614
rect 282306 343378 282542 343614
rect 281986 343058 282222 343294
rect 282306 343058 282542 343294
rect 281986 283378 282222 283614
rect 282306 283378 282542 283614
rect 281986 283058 282222 283294
rect 282306 283058 282542 283294
rect 281986 223378 282222 223614
rect 282306 223378 282542 223614
rect 281986 223058 282222 223294
rect 282306 223058 282542 223294
rect 281986 163378 282222 163614
rect 282306 163378 282542 163614
rect 281986 163058 282222 163294
rect 282306 163058 282542 163294
rect 281986 103378 282222 103614
rect 282306 103378 282542 103614
rect 281986 103058 282222 103294
rect 282306 103058 282542 103294
rect 281986 43378 282222 43614
rect 282306 43378 282542 43614
rect 281986 43058 282222 43294
rect 282306 43058 282542 43294
rect 251986 -6342 252222 -6106
rect 252306 -6342 252542 -6106
rect 251986 -6662 252222 -6426
rect 252306 -6662 252542 -6426
rect 300826 704602 301062 704838
rect 301146 704602 301382 704838
rect 300826 704282 301062 704518
rect 301146 704282 301382 704518
rect 300826 662218 301062 662454
rect 301146 662218 301382 662454
rect 300826 661898 301062 662134
rect 301146 661898 301382 662134
rect 300826 602218 301062 602454
rect 301146 602218 301382 602454
rect 300826 601898 301062 602134
rect 301146 601898 301382 602134
rect 300826 542218 301062 542454
rect 301146 542218 301382 542454
rect 300826 541898 301062 542134
rect 301146 541898 301382 542134
rect 300826 482218 301062 482454
rect 301146 482218 301382 482454
rect 300826 481898 301062 482134
rect 301146 481898 301382 482134
rect 300826 422218 301062 422454
rect 301146 422218 301382 422454
rect 300826 421898 301062 422134
rect 301146 421898 301382 422134
rect 300826 362218 301062 362454
rect 301146 362218 301382 362454
rect 300826 361898 301062 362134
rect 301146 361898 301382 362134
rect 300826 302218 301062 302454
rect 301146 302218 301382 302454
rect 300826 301898 301062 302134
rect 301146 301898 301382 302134
rect 300826 242218 301062 242454
rect 301146 242218 301382 242454
rect 300826 241898 301062 242134
rect 301146 241898 301382 242134
rect 300826 182218 301062 182454
rect 301146 182218 301382 182454
rect 300826 181898 301062 182134
rect 301146 181898 301382 182134
rect 300826 122218 301062 122454
rect 301146 122218 301382 122454
rect 300826 121898 301062 122134
rect 301146 121898 301382 122134
rect 300826 62218 301062 62454
rect 301146 62218 301382 62454
rect 300826 61898 301062 62134
rect 301146 61898 301382 62134
rect 300826 2218 301062 2454
rect 301146 2218 301382 2454
rect 300826 1898 301062 2134
rect 301146 1898 301382 2134
rect 300826 -582 301062 -346
rect 301146 -582 301382 -346
rect 300826 -902 301062 -666
rect 301146 -902 301382 -666
rect 304546 665938 304782 666174
rect 304866 665938 305102 666174
rect 304546 665618 304782 665854
rect 304866 665618 305102 665854
rect 304546 605938 304782 606174
rect 304866 605938 305102 606174
rect 304546 605618 304782 605854
rect 304866 605618 305102 605854
rect 304546 545938 304782 546174
rect 304866 545938 305102 546174
rect 304546 545618 304782 545854
rect 304866 545618 305102 545854
rect 304546 485938 304782 486174
rect 304866 485938 305102 486174
rect 304546 485618 304782 485854
rect 304866 485618 305102 485854
rect 304546 425938 304782 426174
rect 304866 425938 305102 426174
rect 304546 425618 304782 425854
rect 304866 425618 305102 425854
rect 304546 365938 304782 366174
rect 304866 365938 305102 366174
rect 304546 365618 304782 365854
rect 304866 365618 305102 365854
rect 304546 305938 304782 306174
rect 304866 305938 305102 306174
rect 304546 305618 304782 305854
rect 304866 305618 305102 305854
rect 304546 245938 304782 246174
rect 304866 245938 305102 246174
rect 304546 245618 304782 245854
rect 304866 245618 305102 245854
rect 304546 185938 304782 186174
rect 304866 185938 305102 186174
rect 304546 185618 304782 185854
rect 304866 185618 305102 185854
rect 304546 125938 304782 126174
rect 304866 125938 305102 126174
rect 304546 125618 304782 125854
rect 304866 125618 305102 125854
rect 304546 65938 304782 66174
rect 304866 65938 305102 66174
rect 304546 65618 304782 65854
rect 304866 65618 305102 65854
rect 304546 5938 304782 6174
rect 304866 5938 305102 6174
rect 304546 5618 304782 5854
rect 304866 5618 305102 5854
rect 304546 -2502 304782 -2266
rect 304866 -2502 305102 -2266
rect 304546 -2822 304782 -2586
rect 304866 -2822 305102 -2586
rect 308266 669658 308502 669894
rect 308586 669658 308822 669894
rect 308266 669338 308502 669574
rect 308586 669338 308822 669574
rect 308266 609658 308502 609894
rect 308586 609658 308822 609894
rect 308266 609338 308502 609574
rect 308586 609338 308822 609574
rect 308266 549658 308502 549894
rect 308586 549658 308822 549894
rect 308266 549338 308502 549574
rect 308586 549338 308822 549574
rect 308266 489658 308502 489894
rect 308586 489658 308822 489894
rect 308266 489338 308502 489574
rect 308586 489338 308822 489574
rect 308266 429658 308502 429894
rect 308586 429658 308822 429894
rect 308266 429338 308502 429574
rect 308586 429338 308822 429574
rect 308266 369658 308502 369894
rect 308586 369658 308822 369894
rect 308266 369338 308502 369574
rect 308586 369338 308822 369574
rect 308266 309658 308502 309894
rect 308586 309658 308822 309894
rect 308266 309338 308502 309574
rect 308586 309338 308822 309574
rect 308266 249658 308502 249894
rect 308586 249658 308822 249894
rect 308266 249338 308502 249574
rect 308586 249338 308822 249574
rect 308266 189658 308502 189894
rect 308586 189658 308822 189894
rect 308266 189338 308502 189574
rect 308586 189338 308822 189574
rect 308266 129658 308502 129894
rect 308586 129658 308822 129894
rect 308266 129338 308502 129574
rect 308586 129338 308822 129574
rect 308266 69658 308502 69894
rect 308586 69658 308822 69894
rect 308266 69338 308502 69574
rect 308586 69338 308822 69574
rect 308266 9658 308502 9894
rect 308586 9658 308822 9894
rect 308266 9338 308502 9574
rect 308586 9338 308822 9574
rect 308266 -4422 308502 -4186
rect 308586 -4422 308822 -4186
rect 308266 -4742 308502 -4506
rect 308586 -4742 308822 -4506
rect 341986 711322 342222 711558
rect 342306 711322 342542 711558
rect 341986 711002 342222 711238
rect 342306 711002 342542 711238
rect 338266 709402 338502 709638
rect 338586 709402 338822 709638
rect 338266 709082 338502 709318
rect 338586 709082 338822 709318
rect 334546 707482 334782 707718
rect 334866 707482 335102 707718
rect 334546 707162 334782 707398
rect 334866 707162 335102 707398
rect 311986 673378 312222 673614
rect 312306 673378 312542 673614
rect 311986 673058 312222 673294
rect 312306 673058 312542 673294
rect 311986 613378 312222 613614
rect 312306 613378 312542 613614
rect 311986 613058 312222 613294
rect 312306 613058 312542 613294
rect 311986 553378 312222 553614
rect 312306 553378 312542 553614
rect 311986 553058 312222 553294
rect 312306 553058 312542 553294
rect 311986 493378 312222 493614
rect 312306 493378 312542 493614
rect 311986 493058 312222 493294
rect 312306 493058 312542 493294
rect 311986 433378 312222 433614
rect 312306 433378 312542 433614
rect 311986 433058 312222 433294
rect 312306 433058 312542 433294
rect 311986 373378 312222 373614
rect 312306 373378 312542 373614
rect 311986 373058 312222 373294
rect 312306 373058 312542 373294
rect 311986 313378 312222 313614
rect 312306 313378 312542 313614
rect 311986 313058 312222 313294
rect 312306 313058 312542 313294
rect 311986 253378 312222 253614
rect 312306 253378 312542 253614
rect 311986 253058 312222 253294
rect 312306 253058 312542 253294
rect 311986 193378 312222 193614
rect 312306 193378 312542 193614
rect 311986 193058 312222 193294
rect 312306 193058 312542 193294
rect 311986 133378 312222 133614
rect 312306 133378 312542 133614
rect 311986 133058 312222 133294
rect 312306 133058 312542 133294
rect 311986 73378 312222 73614
rect 312306 73378 312542 73614
rect 311986 73058 312222 73294
rect 312306 73058 312542 73294
rect 311986 13378 312222 13614
rect 312306 13378 312542 13614
rect 311986 13058 312222 13294
rect 312306 13058 312542 13294
rect 281986 -7302 282222 -7066
rect 282306 -7302 282542 -7066
rect 281986 -7622 282222 -7386
rect 282306 -7622 282542 -7386
rect 330826 705562 331062 705798
rect 331146 705562 331382 705798
rect 330826 705242 331062 705478
rect 331146 705242 331382 705478
rect 330826 692218 331062 692454
rect 331146 692218 331382 692454
rect 330826 691898 331062 692134
rect 331146 691898 331382 692134
rect 330826 632218 331062 632454
rect 331146 632218 331382 632454
rect 330826 631898 331062 632134
rect 331146 631898 331382 632134
rect 330826 572218 331062 572454
rect 331146 572218 331382 572454
rect 330826 571898 331062 572134
rect 331146 571898 331382 572134
rect 330826 512218 331062 512454
rect 331146 512218 331382 512454
rect 330826 511898 331062 512134
rect 331146 511898 331382 512134
rect 330826 452218 331062 452454
rect 331146 452218 331382 452454
rect 330826 451898 331062 452134
rect 331146 451898 331382 452134
rect 330826 392218 331062 392454
rect 331146 392218 331382 392454
rect 330826 391898 331062 392134
rect 331146 391898 331382 392134
rect 330826 332218 331062 332454
rect 331146 332218 331382 332454
rect 330826 331898 331062 332134
rect 331146 331898 331382 332134
rect 330826 272218 331062 272454
rect 331146 272218 331382 272454
rect 330826 271898 331062 272134
rect 331146 271898 331382 272134
rect 330826 212218 331062 212454
rect 331146 212218 331382 212454
rect 330826 211898 331062 212134
rect 331146 211898 331382 212134
rect 330826 152218 331062 152454
rect 331146 152218 331382 152454
rect 330826 151898 331062 152134
rect 331146 151898 331382 152134
rect 330826 92218 331062 92454
rect 331146 92218 331382 92454
rect 330826 91898 331062 92134
rect 331146 91898 331382 92134
rect 330826 32218 331062 32454
rect 331146 32218 331382 32454
rect 330826 31898 331062 32134
rect 331146 31898 331382 32134
rect 330826 -1542 331062 -1306
rect 331146 -1542 331382 -1306
rect 330826 -1862 331062 -1626
rect 331146 -1862 331382 -1626
rect 334546 695938 334782 696174
rect 334866 695938 335102 696174
rect 334546 695618 334782 695854
rect 334866 695618 335102 695854
rect 334546 635938 334782 636174
rect 334866 635938 335102 636174
rect 334546 635618 334782 635854
rect 334866 635618 335102 635854
rect 334546 575938 334782 576174
rect 334866 575938 335102 576174
rect 334546 575618 334782 575854
rect 334866 575618 335102 575854
rect 334546 515938 334782 516174
rect 334866 515938 335102 516174
rect 334546 515618 334782 515854
rect 334866 515618 335102 515854
rect 334546 455938 334782 456174
rect 334866 455938 335102 456174
rect 334546 455618 334782 455854
rect 334866 455618 335102 455854
rect 334546 395938 334782 396174
rect 334866 395938 335102 396174
rect 334546 395618 334782 395854
rect 334866 395618 335102 395854
rect 334546 335938 334782 336174
rect 334866 335938 335102 336174
rect 334546 335618 334782 335854
rect 334866 335618 335102 335854
rect 334546 275938 334782 276174
rect 334866 275938 335102 276174
rect 334546 275618 334782 275854
rect 334866 275618 335102 275854
rect 334546 215938 334782 216174
rect 334866 215938 335102 216174
rect 334546 215618 334782 215854
rect 334866 215618 335102 215854
rect 334546 155938 334782 156174
rect 334866 155938 335102 156174
rect 334546 155618 334782 155854
rect 334866 155618 335102 155854
rect 334546 95938 334782 96174
rect 334866 95938 335102 96174
rect 334546 95618 334782 95854
rect 334866 95618 335102 95854
rect 334546 35938 334782 36174
rect 334866 35938 335102 36174
rect 334546 35618 334782 35854
rect 334866 35618 335102 35854
rect 334546 -3462 334782 -3226
rect 334866 -3462 335102 -3226
rect 334546 -3782 334782 -3546
rect 334866 -3782 335102 -3546
rect 338266 699658 338502 699894
rect 338586 699658 338822 699894
rect 338266 699338 338502 699574
rect 338586 699338 338822 699574
rect 338266 639658 338502 639894
rect 338586 639658 338822 639894
rect 338266 639338 338502 639574
rect 338586 639338 338822 639574
rect 338266 579658 338502 579894
rect 338586 579658 338822 579894
rect 338266 579338 338502 579574
rect 338586 579338 338822 579574
rect 338266 519658 338502 519894
rect 338586 519658 338822 519894
rect 338266 519338 338502 519574
rect 338586 519338 338822 519574
rect 338266 459658 338502 459894
rect 338586 459658 338822 459894
rect 338266 459338 338502 459574
rect 338586 459338 338822 459574
rect 338266 399658 338502 399894
rect 338586 399658 338822 399894
rect 338266 399338 338502 399574
rect 338586 399338 338822 399574
rect 338266 339658 338502 339894
rect 338586 339658 338822 339894
rect 338266 339338 338502 339574
rect 338586 339338 338822 339574
rect 338266 279658 338502 279894
rect 338586 279658 338822 279894
rect 338266 279338 338502 279574
rect 338586 279338 338822 279574
rect 338266 219658 338502 219894
rect 338586 219658 338822 219894
rect 338266 219338 338502 219574
rect 338586 219338 338822 219574
rect 338266 159658 338502 159894
rect 338586 159658 338822 159894
rect 338266 159338 338502 159574
rect 338586 159338 338822 159574
rect 338266 99658 338502 99894
rect 338586 99658 338822 99894
rect 338266 99338 338502 99574
rect 338586 99338 338822 99574
rect 338266 39658 338502 39894
rect 338586 39658 338822 39894
rect 338266 39338 338502 39574
rect 338586 39338 338822 39574
rect 338266 -5382 338502 -5146
rect 338586 -5382 338822 -5146
rect 338266 -5702 338502 -5466
rect 338586 -5702 338822 -5466
rect 371986 710362 372222 710598
rect 372306 710362 372542 710598
rect 371986 710042 372222 710278
rect 372306 710042 372542 710278
rect 368266 708442 368502 708678
rect 368586 708442 368822 708678
rect 368266 708122 368502 708358
rect 368586 708122 368822 708358
rect 364546 706522 364782 706758
rect 364866 706522 365102 706758
rect 364546 706202 364782 706438
rect 364866 706202 365102 706438
rect 341986 643378 342222 643614
rect 342306 643378 342542 643614
rect 341986 643058 342222 643294
rect 342306 643058 342542 643294
rect 341986 583378 342222 583614
rect 342306 583378 342542 583614
rect 341986 583058 342222 583294
rect 342306 583058 342542 583294
rect 341986 523378 342222 523614
rect 342306 523378 342542 523614
rect 341986 523058 342222 523294
rect 342306 523058 342542 523294
rect 341986 463378 342222 463614
rect 342306 463378 342542 463614
rect 341986 463058 342222 463294
rect 342306 463058 342542 463294
rect 341986 403378 342222 403614
rect 342306 403378 342542 403614
rect 341986 403058 342222 403294
rect 342306 403058 342542 403294
rect 341986 343378 342222 343614
rect 342306 343378 342542 343614
rect 341986 343058 342222 343294
rect 342306 343058 342542 343294
rect 341986 283378 342222 283614
rect 342306 283378 342542 283614
rect 341986 283058 342222 283294
rect 342306 283058 342542 283294
rect 341986 223378 342222 223614
rect 342306 223378 342542 223614
rect 341986 223058 342222 223294
rect 342306 223058 342542 223294
rect 341986 163378 342222 163614
rect 342306 163378 342542 163614
rect 341986 163058 342222 163294
rect 342306 163058 342542 163294
rect 341986 103378 342222 103614
rect 342306 103378 342542 103614
rect 341986 103058 342222 103294
rect 342306 103058 342542 103294
rect 341986 43378 342222 43614
rect 342306 43378 342542 43614
rect 341986 43058 342222 43294
rect 342306 43058 342542 43294
rect 311986 -6342 312222 -6106
rect 312306 -6342 312542 -6106
rect 311986 -6662 312222 -6426
rect 312306 -6662 312542 -6426
rect 360826 704602 361062 704838
rect 361146 704602 361382 704838
rect 360826 704282 361062 704518
rect 361146 704282 361382 704518
rect 360826 662218 361062 662454
rect 361146 662218 361382 662454
rect 360826 661898 361062 662134
rect 361146 661898 361382 662134
rect 360826 602218 361062 602454
rect 361146 602218 361382 602454
rect 360826 601898 361062 602134
rect 361146 601898 361382 602134
rect 360826 542218 361062 542454
rect 361146 542218 361382 542454
rect 360826 541898 361062 542134
rect 361146 541898 361382 542134
rect 360826 482218 361062 482454
rect 361146 482218 361382 482454
rect 360826 481898 361062 482134
rect 361146 481898 361382 482134
rect 360826 422218 361062 422454
rect 361146 422218 361382 422454
rect 360826 421898 361062 422134
rect 361146 421898 361382 422134
rect 360826 362218 361062 362454
rect 361146 362218 361382 362454
rect 360826 361898 361062 362134
rect 361146 361898 361382 362134
rect 360826 302218 361062 302454
rect 361146 302218 361382 302454
rect 360826 301898 361062 302134
rect 361146 301898 361382 302134
rect 360826 242218 361062 242454
rect 361146 242218 361382 242454
rect 360826 241898 361062 242134
rect 361146 241898 361382 242134
rect 360826 182218 361062 182454
rect 361146 182218 361382 182454
rect 360826 181898 361062 182134
rect 361146 181898 361382 182134
rect 360826 122218 361062 122454
rect 361146 122218 361382 122454
rect 360826 121898 361062 122134
rect 361146 121898 361382 122134
rect 360826 62218 361062 62454
rect 361146 62218 361382 62454
rect 360826 61898 361062 62134
rect 361146 61898 361382 62134
rect 360826 2218 361062 2454
rect 361146 2218 361382 2454
rect 360826 1898 361062 2134
rect 361146 1898 361382 2134
rect 360826 -582 361062 -346
rect 361146 -582 361382 -346
rect 360826 -902 361062 -666
rect 361146 -902 361382 -666
rect 364546 665938 364782 666174
rect 364866 665938 365102 666174
rect 364546 665618 364782 665854
rect 364866 665618 365102 665854
rect 364546 605938 364782 606174
rect 364866 605938 365102 606174
rect 364546 605618 364782 605854
rect 364866 605618 365102 605854
rect 364546 545938 364782 546174
rect 364866 545938 365102 546174
rect 364546 545618 364782 545854
rect 364866 545618 365102 545854
rect 364546 485938 364782 486174
rect 364866 485938 365102 486174
rect 364546 485618 364782 485854
rect 364866 485618 365102 485854
rect 364546 425938 364782 426174
rect 364866 425938 365102 426174
rect 364546 425618 364782 425854
rect 364866 425618 365102 425854
rect 364546 365938 364782 366174
rect 364866 365938 365102 366174
rect 364546 365618 364782 365854
rect 364866 365618 365102 365854
rect 364546 305938 364782 306174
rect 364866 305938 365102 306174
rect 364546 305618 364782 305854
rect 364866 305618 365102 305854
rect 364546 245938 364782 246174
rect 364866 245938 365102 246174
rect 364546 245618 364782 245854
rect 364866 245618 365102 245854
rect 364546 185938 364782 186174
rect 364866 185938 365102 186174
rect 364546 185618 364782 185854
rect 364866 185618 365102 185854
rect 364546 125938 364782 126174
rect 364866 125938 365102 126174
rect 364546 125618 364782 125854
rect 364866 125618 365102 125854
rect 364546 65938 364782 66174
rect 364866 65938 365102 66174
rect 364546 65618 364782 65854
rect 364866 65618 365102 65854
rect 364546 5938 364782 6174
rect 364866 5938 365102 6174
rect 364546 5618 364782 5854
rect 364866 5618 365102 5854
rect 364546 -2502 364782 -2266
rect 364866 -2502 365102 -2266
rect 364546 -2822 364782 -2586
rect 364866 -2822 365102 -2586
rect 368266 669658 368502 669894
rect 368586 669658 368822 669894
rect 368266 669338 368502 669574
rect 368586 669338 368822 669574
rect 368266 609658 368502 609894
rect 368586 609658 368822 609894
rect 368266 609338 368502 609574
rect 368586 609338 368822 609574
rect 368266 549658 368502 549894
rect 368586 549658 368822 549894
rect 368266 549338 368502 549574
rect 368586 549338 368822 549574
rect 368266 489658 368502 489894
rect 368586 489658 368822 489894
rect 368266 489338 368502 489574
rect 368586 489338 368822 489574
rect 368266 429658 368502 429894
rect 368586 429658 368822 429894
rect 368266 429338 368502 429574
rect 368586 429338 368822 429574
rect 368266 369658 368502 369894
rect 368586 369658 368822 369894
rect 368266 369338 368502 369574
rect 368586 369338 368822 369574
rect 368266 309658 368502 309894
rect 368586 309658 368822 309894
rect 368266 309338 368502 309574
rect 368586 309338 368822 309574
rect 368266 249658 368502 249894
rect 368586 249658 368822 249894
rect 368266 249338 368502 249574
rect 368586 249338 368822 249574
rect 368266 189658 368502 189894
rect 368586 189658 368822 189894
rect 368266 189338 368502 189574
rect 368586 189338 368822 189574
rect 368266 129658 368502 129894
rect 368586 129658 368822 129894
rect 368266 129338 368502 129574
rect 368586 129338 368822 129574
rect 368266 69658 368502 69894
rect 368586 69658 368822 69894
rect 368266 69338 368502 69574
rect 368586 69338 368822 69574
rect 368266 9658 368502 9894
rect 368586 9658 368822 9894
rect 368266 9338 368502 9574
rect 368586 9338 368822 9574
rect 368266 -4422 368502 -4186
rect 368586 -4422 368822 -4186
rect 368266 -4742 368502 -4506
rect 368586 -4742 368822 -4506
rect 401986 711322 402222 711558
rect 402306 711322 402542 711558
rect 401986 711002 402222 711238
rect 402306 711002 402542 711238
rect 398266 709402 398502 709638
rect 398586 709402 398822 709638
rect 398266 709082 398502 709318
rect 398586 709082 398822 709318
rect 394546 707482 394782 707718
rect 394866 707482 395102 707718
rect 394546 707162 394782 707398
rect 394866 707162 395102 707398
rect 371986 673378 372222 673614
rect 372306 673378 372542 673614
rect 371986 673058 372222 673294
rect 372306 673058 372542 673294
rect 371986 613378 372222 613614
rect 372306 613378 372542 613614
rect 371986 613058 372222 613294
rect 372306 613058 372542 613294
rect 371986 553378 372222 553614
rect 372306 553378 372542 553614
rect 371986 553058 372222 553294
rect 372306 553058 372542 553294
rect 371986 493378 372222 493614
rect 372306 493378 372542 493614
rect 371986 493058 372222 493294
rect 372306 493058 372542 493294
rect 371986 433378 372222 433614
rect 372306 433378 372542 433614
rect 371986 433058 372222 433294
rect 372306 433058 372542 433294
rect 371986 373378 372222 373614
rect 372306 373378 372542 373614
rect 371986 373058 372222 373294
rect 372306 373058 372542 373294
rect 371986 313378 372222 313614
rect 372306 313378 372542 313614
rect 371986 313058 372222 313294
rect 372306 313058 372542 313294
rect 371986 253378 372222 253614
rect 372306 253378 372542 253614
rect 371986 253058 372222 253294
rect 372306 253058 372542 253294
rect 371986 193378 372222 193614
rect 372306 193378 372542 193614
rect 371986 193058 372222 193294
rect 372306 193058 372542 193294
rect 371986 133378 372222 133614
rect 372306 133378 372542 133614
rect 371986 133058 372222 133294
rect 372306 133058 372542 133294
rect 371986 73378 372222 73614
rect 372306 73378 372542 73614
rect 371986 73058 372222 73294
rect 372306 73058 372542 73294
rect 371986 13378 372222 13614
rect 372306 13378 372542 13614
rect 371986 13058 372222 13294
rect 372306 13058 372542 13294
rect 341986 -7302 342222 -7066
rect 342306 -7302 342542 -7066
rect 341986 -7622 342222 -7386
rect 342306 -7622 342542 -7386
rect 390826 705562 391062 705798
rect 391146 705562 391382 705798
rect 390826 705242 391062 705478
rect 391146 705242 391382 705478
rect 390826 692218 391062 692454
rect 391146 692218 391382 692454
rect 390826 691898 391062 692134
rect 391146 691898 391382 692134
rect 390826 632218 391062 632454
rect 391146 632218 391382 632454
rect 390826 631898 391062 632134
rect 391146 631898 391382 632134
rect 390826 572218 391062 572454
rect 391146 572218 391382 572454
rect 390826 571898 391062 572134
rect 391146 571898 391382 572134
rect 390826 512218 391062 512454
rect 391146 512218 391382 512454
rect 390826 511898 391062 512134
rect 391146 511898 391382 512134
rect 390826 452218 391062 452454
rect 391146 452218 391382 452454
rect 390826 451898 391062 452134
rect 391146 451898 391382 452134
rect 390826 392218 391062 392454
rect 391146 392218 391382 392454
rect 390826 391898 391062 392134
rect 391146 391898 391382 392134
rect 390826 332218 391062 332454
rect 391146 332218 391382 332454
rect 390826 331898 391062 332134
rect 391146 331898 391382 332134
rect 390826 272218 391062 272454
rect 391146 272218 391382 272454
rect 390826 271898 391062 272134
rect 391146 271898 391382 272134
rect 390826 212218 391062 212454
rect 391146 212218 391382 212454
rect 390826 211898 391062 212134
rect 391146 211898 391382 212134
rect 390826 152218 391062 152454
rect 391146 152218 391382 152454
rect 390826 151898 391062 152134
rect 391146 151898 391382 152134
rect 390826 92218 391062 92454
rect 391146 92218 391382 92454
rect 390826 91898 391062 92134
rect 391146 91898 391382 92134
rect 390826 32218 391062 32454
rect 391146 32218 391382 32454
rect 390826 31898 391062 32134
rect 391146 31898 391382 32134
rect 390826 -1542 391062 -1306
rect 391146 -1542 391382 -1306
rect 390826 -1862 391062 -1626
rect 391146 -1862 391382 -1626
rect 394546 695938 394782 696174
rect 394866 695938 395102 696174
rect 394546 695618 394782 695854
rect 394866 695618 395102 695854
rect 394546 635938 394782 636174
rect 394866 635938 395102 636174
rect 394546 635618 394782 635854
rect 394866 635618 395102 635854
rect 394546 575938 394782 576174
rect 394866 575938 395102 576174
rect 394546 575618 394782 575854
rect 394866 575618 395102 575854
rect 394546 515938 394782 516174
rect 394866 515938 395102 516174
rect 394546 515618 394782 515854
rect 394866 515618 395102 515854
rect 394546 455938 394782 456174
rect 394866 455938 395102 456174
rect 394546 455618 394782 455854
rect 394866 455618 395102 455854
rect 394546 395938 394782 396174
rect 394866 395938 395102 396174
rect 394546 395618 394782 395854
rect 394866 395618 395102 395854
rect 394546 335938 394782 336174
rect 394866 335938 395102 336174
rect 394546 335618 394782 335854
rect 394866 335618 395102 335854
rect 394546 275938 394782 276174
rect 394866 275938 395102 276174
rect 394546 275618 394782 275854
rect 394866 275618 395102 275854
rect 394546 215938 394782 216174
rect 394866 215938 395102 216174
rect 394546 215618 394782 215854
rect 394866 215618 395102 215854
rect 394546 155938 394782 156174
rect 394866 155938 395102 156174
rect 394546 155618 394782 155854
rect 394866 155618 395102 155854
rect 394546 95938 394782 96174
rect 394866 95938 395102 96174
rect 394546 95618 394782 95854
rect 394866 95618 395102 95854
rect 394546 35938 394782 36174
rect 394866 35938 395102 36174
rect 394546 35618 394782 35854
rect 394866 35618 395102 35854
rect 394546 -3462 394782 -3226
rect 394866 -3462 395102 -3226
rect 394546 -3782 394782 -3546
rect 394866 -3782 395102 -3546
rect 398266 699658 398502 699894
rect 398586 699658 398822 699894
rect 398266 699338 398502 699574
rect 398586 699338 398822 699574
rect 398266 639658 398502 639894
rect 398586 639658 398822 639894
rect 398266 639338 398502 639574
rect 398586 639338 398822 639574
rect 398266 579658 398502 579894
rect 398586 579658 398822 579894
rect 398266 579338 398502 579574
rect 398586 579338 398822 579574
rect 398266 519658 398502 519894
rect 398586 519658 398822 519894
rect 398266 519338 398502 519574
rect 398586 519338 398822 519574
rect 398266 459658 398502 459894
rect 398586 459658 398822 459894
rect 398266 459338 398502 459574
rect 398586 459338 398822 459574
rect 398266 399658 398502 399894
rect 398586 399658 398822 399894
rect 398266 399338 398502 399574
rect 398586 399338 398822 399574
rect 398266 339658 398502 339894
rect 398586 339658 398822 339894
rect 398266 339338 398502 339574
rect 398586 339338 398822 339574
rect 398266 279658 398502 279894
rect 398586 279658 398822 279894
rect 398266 279338 398502 279574
rect 398586 279338 398822 279574
rect 398266 219658 398502 219894
rect 398586 219658 398822 219894
rect 398266 219338 398502 219574
rect 398586 219338 398822 219574
rect 398266 159658 398502 159894
rect 398586 159658 398822 159894
rect 398266 159338 398502 159574
rect 398586 159338 398822 159574
rect 398266 99658 398502 99894
rect 398586 99658 398822 99894
rect 398266 99338 398502 99574
rect 398586 99338 398822 99574
rect 398266 39658 398502 39894
rect 398586 39658 398822 39894
rect 398266 39338 398502 39574
rect 398586 39338 398822 39574
rect 398266 -5382 398502 -5146
rect 398586 -5382 398822 -5146
rect 398266 -5702 398502 -5466
rect 398586 -5702 398822 -5466
rect 431986 710362 432222 710598
rect 432306 710362 432542 710598
rect 431986 710042 432222 710278
rect 432306 710042 432542 710278
rect 428266 708442 428502 708678
rect 428586 708442 428822 708678
rect 428266 708122 428502 708358
rect 428586 708122 428822 708358
rect 424546 706522 424782 706758
rect 424866 706522 425102 706758
rect 424546 706202 424782 706438
rect 424866 706202 425102 706438
rect 401986 643378 402222 643614
rect 402306 643378 402542 643614
rect 401986 643058 402222 643294
rect 402306 643058 402542 643294
rect 401986 583378 402222 583614
rect 402306 583378 402542 583614
rect 401986 583058 402222 583294
rect 402306 583058 402542 583294
rect 401986 523378 402222 523614
rect 402306 523378 402542 523614
rect 401986 523058 402222 523294
rect 402306 523058 402542 523294
rect 401986 463378 402222 463614
rect 402306 463378 402542 463614
rect 401986 463058 402222 463294
rect 402306 463058 402542 463294
rect 401986 403378 402222 403614
rect 402306 403378 402542 403614
rect 401986 403058 402222 403294
rect 402306 403058 402542 403294
rect 401986 343378 402222 343614
rect 402306 343378 402542 343614
rect 401986 343058 402222 343294
rect 402306 343058 402542 343294
rect 401986 283378 402222 283614
rect 402306 283378 402542 283614
rect 401986 283058 402222 283294
rect 402306 283058 402542 283294
rect 401986 223378 402222 223614
rect 402306 223378 402542 223614
rect 401986 223058 402222 223294
rect 402306 223058 402542 223294
rect 401986 163378 402222 163614
rect 402306 163378 402542 163614
rect 401986 163058 402222 163294
rect 402306 163058 402542 163294
rect 401986 103378 402222 103614
rect 402306 103378 402542 103614
rect 401986 103058 402222 103294
rect 402306 103058 402542 103294
rect 401986 43378 402222 43614
rect 402306 43378 402542 43614
rect 401986 43058 402222 43294
rect 402306 43058 402542 43294
rect 371986 -6342 372222 -6106
rect 372306 -6342 372542 -6106
rect 371986 -6662 372222 -6426
rect 372306 -6662 372542 -6426
rect 420826 704602 421062 704838
rect 421146 704602 421382 704838
rect 420826 704282 421062 704518
rect 421146 704282 421382 704518
rect 420826 662218 421062 662454
rect 421146 662218 421382 662454
rect 420826 661898 421062 662134
rect 421146 661898 421382 662134
rect 420826 602218 421062 602454
rect 421146 602218 421382 602454
rect 420826 601898 421062 602134
rect 421146 601898 421382 602134
rect 420826 542218 421062 542454
rect 421146 542218 421382 542454
rect 420826 541898 421062 542134
rect 421146 541898 421382 542134
rect 420826 482218 421062 482454
rect 421146 482218 421382 482454
rect 420826 481898 421062 482134
rect 421146 481898 421382 482134
rect 420826 422218 421062 422454
rect 421146 422218 421382 422454
rect 420826 421898 421062 422134
rect 421146 421898 421382 422134
rect 420826 362218 421062 362454
rect 421146 362218 421382 362454
rect 420826 361898 421062 362134
rect 421146 361898 421382 362134
rect 420826 302218 421062 302454
rect 421146 302218 421382 302454
rect 420826 301898 421062 302134
rect 421146 301898 421382 302134
rect 420826 242218 421062 242454
rect 421146 242218 421382 242454
rect 420826 241898 421062 242134
rect 421146 241898 421382 242134
rect 420826 182218 421062 182454
rect 421146 182218 421382 182454
rect 420826 181898 421062 182134
rect 421146 181898 421382 182134
rect 420826 122218 421062 122454
rect 421146 122218 421382 122454
rect 420826 121898 421062 122134
rect 421146 121898 421382 122134
rect 420826 62218 421062 62454
rect 421146 62218 421382 62454
rect 420826 61898 421062 62134
rect 421146 61898 421382 62134
rect 420826 2218 421062 2454
rect 421146 2218 421382 2454
rect 420826 1898 421062 2134
rect 421146 1898 421382 2134
rect 420826 -582 421062 -346
rect 421146 -582 421382 -346
rect 420826 -902 421062 -666
rect 421146 -902 421382 -666
rect 424546 665938 424782 666174
rect 424866 665938 425102 666174
rect 424546 665618 424782 665854
rect 424866 665618 425102 665854
rect 424546 605938 424782 606174
rect 424866 605938 425102 606174
rect 424546 605618 424782 605854
rect 424866 605618 425102 605854
rect 424546 545938 424782 546174
rect 424866 545938 425102 546174
rect 424546 545618 424782 545854
rect 424866 545618 425102 545854
rect 424546 485938 424782 486174
rect 424866 485938 425102 486174
rect 424546 485618 424782 485854
rect 424866 485618 425102 485854
rect 424546 425938 424782 426174
rect 424866 425938 425102 426174
rect 424546 425618 424782 425854
rect 424866 425618 425102 425854
rect 424546 365938 424782 366174
rect 424866 365938 425102 366174
rect 424546 365618 424782 365854
rect 424866 365618 425102 365854
rect 424546 305938 424782 306174
rect 424866 305938 425102 306174
rect 424546 305618 424782 305854
rect 424866 305618 425102 305854
rect 424546 245938 424782 246174
rect 424866 245938 425102 246174
rect 424546 245618 424782 245854
rect 424866 245618 425102 245854
rect 424546 185938 424782 186174
rect 424866 185938 425102 186174
rect 424546 185618 424782 185854
rect 424866 185618 425102 185854
rect 424546 125938 424782 126174
rect 424866 125938 425102 126174
rect 424546 125618 424782 125854
rect 424866 125618 425102 125854
rect 424546 65938 424782 66174
rect 424866 65938 425102 66174
rect 424546 65618 424782 65854
rect 424866 65618 425102 65854
rect 424546 5938 424782 6174
rect 424866 5938 425102 6174
rect 424546 5618 424782 5854
rect 424866 5618 425102 5854
rect 424546 -2502 424782 -2266
rect 424866 -2502 425102 -2266
rect 424546 -2822 424782 -2586
rect 424866 -2822 425102 -2586
rect 428266 669658 428502 669894
rect 428586 669658 428822 669894
rect 428266 669338 428502 669574
rect 428586 669338 428822 669574
rect 428266 609658 428502 609894
rect 428586 609658 428822 609894
rect 428266 609338 428502 609574
rect 428586 609338 428822 609574
rect 428266 549658 428502 549894
rect 428586 549658 428822 549894
rect 428266 549338 428502 549574
rect 428586 549338 428822 549574
rect 428266 489658 428502 489894
rect 428586 489658 428822 489894
rect 428266 489338 428502 489574
rect 428586 489338 428822 489574
rect 428266 429658 428502 429894
rect 428586 429658 428822 429894
rect 428266 429338 428502 429574
rect 428586 429338 428822 429574
rect 428266 369658 428502 369894
rect 428586 369658 428822 369894
rect 428266 369338 428502 369574
rect 428586 369338 428822 369574
rect 428266 309658 428502 309894
rect 428586 309658 428822 309894
rect 428266 309338 428502 309574
rect 428586 309338 428822 309574
rect 428266 249658 428502 249894
rect 428586 249658 428822 249894
rect 428266 249338 428502 249574
rect 428586 249338 428822 249574
rect 428266 189658 428502 189894
rect 428586 189658 428822 189894
rect 428266 189338 428502 189574
rect 428586 189338 428822 189574
rect 428266 129658 428502 129894
rect 428586 129658 428822 129894
rect 428266 129338 428502 129574
rect 428586 129338 428822 129574
rect 428266 69658 428502 69894
rect 428586 69658 428822 69894
rect 428266 69338 428502 69574
rect 428586 69338 428822 69574
rect 428266 9658 428502 9894
rect 428586 9658 428822 9894
rect 428266 9338 428502 9574
rect 428586 9338 428822 9574
rect 428266 -4422 428502 -4186
rect 428586 -4422 428822 -4186
rect 428266 -4742 428502 -4506
rect 428586 -4742 428822 -4506
rect 461986 711322 462222 711558
rect 462306 711322 462542 711558
rect 461986 711002 462222 711238
rect 462306 711002 462542 711238
rect 458266 709402 458502 709638
rect 458586 709402 458822 709638
rect 458266 709082 458502 709318
rect 458586 709082 458822 709318
rect 454546 707482 454782 707718
rect 454866 707482 455102 707718
rect 454546 707162 454782 707398
rect 454866 707162 455102 707398
rect 431986 673378 432222 673614
rect 432306 673378 432542 673614
rect 431986 673058 432222 673294
rect 432306 673058 432542 673294
rect 431986 613378 432222 613614
rect 432306 613378 432542 613614
rect 431986 613058 432222 613294
rect 432306 613058 432542 613294
rect 431986 553378 432222 553614
rect 432306 553378 432542 553614
rect 431986 553058 432222 553294
rect 432306 553058 432542 553294
rect 431986 493378 432222 493614
rect 432306 493378 432542 493614
rect 431986 493058 432222 493294
rect 432306 493058 432542 493294
rect 431986 433378 432222 433614
rect 432306 433378 432542 433614
rect 431986 433058 432222 433294
rect 432306 433058 432542 433294
rect 431986 373378 432222 373614
rect 432306 373378 432542 373614
rect 431986 373058 432222 373294
rect 432306 373058 432542 373294
rect 431986 313378 432222 313614
rect 432306 313378 432542 313614
rect 431986 313058 432222 313294
rect 432306 313058 432542 313294
rect 431986 253378 432222 253614
rect 432306 253378 432542 253614
rect 431986 253058 432222 253294
rect 432306 253058 432542 253294
rect 431986 193378 432222 193614
rect 432306 193378 432542 193614
rect 431986 193058 432222 193294
rect 432306 193058 432542 193294
rect 431986 133378 432222 133614
rect 432306 133378 432542 133614
rect 431986 133058 432222 133294
rect 432306 133058 432542 133294
rect 431986 73378 432222 73614
rect 432306 73378 432542 73614
rect 431986 73058 432222 73294
rect 432306 73058 432542 73294
rect 431986 13378 432222 13614
rect 432306 13378 432542 13614
rect 431986 13058 432222 13294
rect 432306 13058 432542 13294
rect 401986 -7302 402222 -7066
rect 402306 -7302 402542 -7066
rect 401986 -7622 402222 -7386
rect 402306 -7622 402542 -7386
rect 450826 705562 451062 705798
rect 451146 705562 451382 705798
rect 450826 705242 451062 705478
rect 451146 705242 451382 705478
rect 450826 692218 451062 692454
rect 451146 692218 451382 692454
rect 450826 691898 451062 692134
rect 451146 691898 451382 692134
rect 450826 632218 451062 632454
rect 451146 632218 451382 632454
rect 450826 631898 451062 632134
rect 451146 631898 451382 632134
rect 450826 572218 451062 572454
rect 451146 572218 451382 572454
rect 450826 571898 451062 572134
rect 451146 571898 451382 572134
rect 450826 512218 451062 512454
rect 451146 512218 451382 512454
rect 450826 511898 451062 512134
rect 451146 511898 451382 512134
rect 450826 452218 451062 452454
rect 451146 452218 451382 452454
rect 450826 451898 451062 452134
rect 451146 451898 451382 452134
rect 450826 392218 451062 392454
rect 451146 392218 451382 392454
rect 450826 391898 451062 392134
rect 451146 391898 451382 392134
rect 450826 332218 451062 332454
rect 451146 332218 451382 332454
rect 450826 331898 451062 332134
rect 451146 331898 451382 332134
rect 450826 272218 451062 272454
rect 451146 272218 451382 272454
rect 450826 271898 451062 272134
rect 451146 271898 451382 272134
rect 450826 212218 451062 212454
rect 451146 212218 451382 212454
rect 450826 211898 451062 212134
rect 451146 211898 451382 212134
rect 450826 152218 451062 152454
rect 451146 152218 451382 152454
rect 450826 151898 451062 152134
rect 451146 151898 451382 152134
rect 450826 92218 451062 92454
rect 451146 92218 451382 92454
rect 450826 91898 451062 92134
rect 451146 91898 451382 92134
rect 450826 32218 451062 32454
rect 451146 32218 451382 32454
rect 450826 31898 451062 32134
rect 451146 31898 451382 32134
rect 450826 -1542 451062 -1306
rect 451146 -1542 451382 -1306
rect 450826 -1862 451062 -1626
rect 451146 -1862 451382 -1626
rect 454546 695938 454782 696174
rect 454866 695938 455102 696174
rect 454546 695618 454782 695854
rect 454866 695618 455102 695854
rect 454546 635938 454782 636174
rect 454866 635938 455102 636174
rect 454546 635618 454782 635854
rect 454866 635618 455102 635854
rect 454546 575938 454782 576174
rect 454866 575938 455102 576174
rect 454546 575618 454782 575854
rect 454866 575618 455102 575854
rect 454546 515938 454782 516174
rect 454866 515938 455102 516174
rect 454546 515618 454782 515854
rect 454866 515618 455102 515854
rect 454546 455938 454782 456174
rect 454866 455938 455102 456174
rect 454546 455618 454782 455854
rect 454866 455618 455102 455854
rect 454546 395938 454782 396174
rect 454866 395938 455102 396174
rect 454546 395618 454782 395854
rect 454866 395618 455102 395854
rect 454546 335938 454782 336174
rect 454866 335938 455102 336174
rect 454546 335618 454782 335854
rect 454866 335618 455102 335854
rect 454546 275938 454782 276174
rect 454866 275938 455102 276174
rect 454546 275618 454782 275854
rect 454866 275618 455102 275854
rect 454546 215938 454782 216174
rect 454866 215938 455102 216174
rect 454546 215618 454782 215854
rect 454866 215618 455102 215854
rect 454546 155938 454782 156174
rect 454866 155938 455102 156174
rect 454546 155618 454782 155854
rect 454866 155618 455102 155854
rect 454546 95938 454782 96174
rect 454866 95938 455102 96174
rect 454546 95618 454782 95854
rect 454866 95618 455102 95854
rect 454546 35938 454782 36174
rect 454866 35938 455102 36174
rect 454546 35618 454782 35854
rect 454866 35618 455102 35854
rect 454546 -3462 454782 -3226
rect 454866 -3462 455102 -3226
rect 454546 -3782 454782 -3546
rect 454866 -3782 455102 -3546
rect 458266 699658 458502 699894
rect 458586 699658 458822 699894
rect 458266 699338 458502 699574
rect 458586 699338 458822 699574
rect 458266 639658 458502 639894
rect 458586 639658 458822 639894
rect 458266 639338 458502 639574
rect 458586 639338 458822 639574
rect 458266 579658 458502 579894
rect 458586 579658 458822 579894
rect 458266 579338 458502 579574
rect 458586 579338 458822 579574
rect 458266 519658 458502 519894
rect 458586 519658 458822 519894
rect 458266 519338 458502 519574
rect 458586 519338 458822 519574
rect 458266 459658 458502 459894
rect 458586 459658 458822 459894
rect 458266 459338 458502 459574
rect 458586 459338 458822 459574
rect 458266 399658 458502 399894
rect 458586 399658 458822 399894
rect 458266 399338 458502 399574
rect 458586 399338 458822 399574
rect 458266 339658 458502 339894
rect 458586 339658 458822 339894
rect 458266 339338 458502 339574
rect 458586 339338 458822 339574
rect 458266 279658 458502 279894
rect 458586 279658 458822 279894
rect 458266 279338 458502 279574
rect 458586 279338 458822 279574
rect 458266 219658 458502 219894
rect 458586 219658 458822 219894
rect 458266 219338 458502 219574
rect 458586 219338 458822 219574
rect 458266 159658 458502 159894
rect 458586 159658 458822 159894
rect 458266 159338 458502 159574
rect 458586 159338 458822 159574
rect 458266 99658 458502 99894
rect 458586 99658 458822 99894
rect 458266 99338 458502 99574
rect 458586 99338 458822 99574
rect 458266 39658 458502 39894
rect 458586 39658 458822 39894
rect 458266 39338 458502 39574
rect 458586 39338 458822 39574
rect 458266 -5382 458502 -5146
rect 458586 -5382 458822 -5146
rect 458266 -5702 458502 -5466
rect 458586 -5702 458822 -5466
rect 491986 710362 492222 710598
rect 492306 710362 492542 710598
rect 491986 710042 492222 710278
rect 492306 710042 492542 710278
rect 488266 708442 488502 708678
rect 488586 708442 488822 708678
rect 488266 708122 488502 708358
rect 488586 708122 488822 708358
rect 484546 706522 484782 706758
rect 484866 706522 485102 706758
rect 484546 706202 484782 706438
rect 484866 706202 485102 706438
rect 461986 643378 462222 643614
rect 462306 643378 462542 643614
rect 461986 643058 462222 643294
rect 462306 643058 462542 643294
rect 461986 583378 462222 583614
rect 462306 583378 462542 583614
rect 461986 583058 462222 583294
rect 462306 583058 462542 583294
rect 461986 523378 462222 523614
rect 462306 523378 462542 523614
rect 461986 523058 462222 523294
rect 462306 523058 462542 523294
rect 461986 463378 462222 463614
rect 462306 463378 462542 463614
rect 461986 463058 462222 463294
rect 462306 463058 462542 463294
rect 461986 403378 462222 403614
rect 462306 403378 462542 403614
rect 461986 403058 462222 403294
rect 462306 403058 462542 403294
rect 461986 343378 462222 343614
rect 462306 343378 462542 343614
rect 461986 343058 462222 343294
rect 462306 343058 462542 343294
rect 461986 283378 462222 283614
rect 462306 283378 462542 283614
rect 461986 283058 462222 283294
rect 462306 283058 462542 283294
rect 461986 223378 462222 223614
rect 462306 223378 462542 223614
rect 461986 223058 462222 223294
rect 462306 223058 462542 223294
rect 461986 163378 462222 163614
rect 462306 163378 462542 163614
rect 461986 163058 462222 163294
rect 462306 163058 462542 163294
rect 461986 103378 462222 103614
rect 462306 103378 462542 103614
rect 461986 103058 462222 103294
rect 462306 103058 462542 103294
rect 461986 43378 462222 43614
rect 462306 43378 462542 43614
rect 461986 43058 462222 43294
rect 462306 43058 462542 43294
rect 431986 -6342 432222 -6106
rect 432306 -6342 432542 -6106
rect 431986 -6662 432222 -6426
rect 432306 -6662 432542 -6426
rect 480826 704602 481062 704838
rect 481146 704602 481382 704838
rect 480826 704282 481062 704518
rect 481146 704282 481382 704518
rect 480826 662218 481062 662454
rect 481146 662218 481382 662454
rect 480826 661898 481062 662134
rect 481146 661898 481382 662134
rect 480826 602218 481062 602454
rect 481146 602218 481382 602454
rect 480826 601898 481062 602134
rect 481146 601898 481382 602134
rect 480826 542218 481062 542454
rect 481146 542218 481382 542454
rect 480826 541898 481062 542134
rect 481146 541898 481382 542134
rect 480826 482218 481062 482454
rect 481146 482218 481382 482454
rect 480826 481898 481062 482134
rect 481146 481898 481382 482134
rect 480826 422218 481062 422454
rect 481146 422218 481382 422454
rect 480826 421898 481062 422134
rect 481146 421898 481382 422134
rect 480826 362218 481062 362454
rect 481146 362218 481382 362454
rect 480826 361898 481062 362134
rect 481146 361898 481382 362134
rect 480826 302218 481062 302454
rect 481146 302218 481382 302454
rect 480826 301898 481062 302134
rect 481146 301898 481382 302134
rect 480826 242218 481062 242454
rect 481146 242218 481382 242454
rect 480826 241898 481062 242134
rect 481146 241898 481382 242134
rect 480826 182218 481062 182454
rect 481146 182218 481382 182454
rect 480826 181898 481062 182134
rect 481146 181898 481382 182134
rect 480826 122218 481062 122454
rect 481146 122218 481382 122454
rect 480826 121898 481062 122134
rect 481146 121898 481382 122134
rect 480826 62218 481062 62454
rect 481146 62218 481382 62454
rect 480826 61898 481062 62134
rect 481146 61898 481382 62134
rect 480826 2218 481062 2454
rect 481146 2218 481382 2454
rect 480826 1898 481062 2134
rect 481146 1898 481382 2134
rect 480826 -582 481062 -346
rect 481146 -582 481382 -346
rect 480826 -902 481062 -666
rect 481146 -902 481382 -666
rect 484546 665938 484782 666174
rect 484866 665938 485102 666174
rect 484546 665618 484782 665854
rect 484866 665618 485102 665854
rect 484546 605938 484782 606174
rect 484866 605938 485102 606174
rect 484546 605618 484782 605854
rect 484866 605618 485102 605854
rect 484546 545938 484782 546174
rect 484866 545938 485102 546174
rect 484546 545618 484782 545854
rect 484866 545618 485102 545854
rect 484546 485938 484782 486174
rect 484866 485938 485102 486174
rect 484546 485618 484782 485854
rect 484866 485618 485102 485854
rect 484546 425938 484782 426174
rect 484866 425938 485102 426174
rect 484546 425618 484782 425854
rect 484866 425618 485102 425854
rect 484546 365938 484782 366174
rect 484866 365938 485102 366174
rect 484546 365618 484782 365854
rect 484866 365618 485102 365854
rect 484546 305938 484782 306174
rect 484866 305938 485102 306174
rect 484546 305618 484782 305854
rect 484866 305618 485102 305854
rect 484546 245938 484782 246174
rect 484866 245938 485102 246174
rect 484546 245618 484782 245854
rect 484866 245618 485102 245854
rect 484546 185938 484782 186174
rect 484866 185938 485102 186174
rect 484546 185618 484782 185854
rect 484866 185618 485102 185854
rect 484546 125938 484782 126174
rect 484866 125938 485102 126174
rect 484546 125618 484782 125854
rect 484866 125618 485102 125854
rect 484546 65938 484782 66174
rect 484866 65938 485102 66174
rect 484546 65618 484782 65854
rect 484866 65618 485102 65854
rect 484546 5938 484782 6174
rect 484866 5938 485102 6174
rect 484546 5618 484782 5854
rect 484866 5618 485102 5854
rect 484546 -2502 484782 -2266
rect 484866 -2502 485102 -2266
rect 484546 -2822 484782 -2586
rect 484866 -2822 485102 -2586
rect 488266 669658 488502 669894
rect 488586 669658 488822 669894
rect 488266 669338 488502 669574
rect 488586 669338 488822 669574
rect 488266 609658 488502 609894
rect 488586 609658 488822 609894
rect 488266 609338 488502 609574
rect 488586 609338 488822 609574
rect 488266 549658 488502 549894
rect 488586 549658 488822 549894
rect 488266 549338 488502 549574
rect 488586 549338 488822 549574
rect 488266 489658 488502 489894
rect 488586 489658 488822 489894
rect 488266 489338 488502 489574
rect 488586 489338 488822 489574
rect 488266 429658 488502 429894
rect 488586 429658 488822 429894
rect 488266 429338 488502 429574
rect 488586 429338 488822 429574
rect 488266 369658 488502 369894
rect 488586 369658 488822 369894
rect 488266 369338 488502 369574
rect 488586 369338 488822 369574
rect 488266 309658 488502 309894
rect 488586 309658 488822 309894
rect 488266 309338 488502 309574
rect 488586 309338 488822 309574
rect 488266 249658 488502 249894
rect 488586 249658 488822 249894
rect 488266 249338 488502 249574
rect 488586 249338 488822 249574
rect 488266 189658 488502 189894
rect 488586 189658 488822 189894
rect 488266 189338 488502 189574
rect 488586 189338 488822 189574
rect 488266 129658 488502 129894
rect 488586 129658 488822 129894
rect 488266 129338 488502 129574
rect 488586 129338 488822 129574
rect 488266 69658 488502 69894
rect 488586 69658 488822 69894
rect 488266 69338 488502 69574
rect 488586 69338 488822 69574
rect 488266 9658 488502 9894
rect 488586 9658 488822 9894
rect 488266 9338 488502 9574
rect 488586 9338 488822 9574
rect 488266 -4422 488502 -4186
rect 488586 -4422 488822 -4186
rect 488266 -4742 488502 -4506
rect 488586 -4742 488822 -4506
rect 521986 711322 522222 711558
rect 522306 711322 522542 711558
rect 521986 711002 522222 711238
rect 522306 711002 522542 711238
rect 518266 709402 518502 709638
rect 518586 709402 518822 709638
rect 518266 709082 518502 709318
rect 518586 709082 518822 709318
rect 514546 707482 514782 707718
rect 514866 707482 515102 707718
rect 514546 707162 514782 707398
rect 514866 707162 515102 707398
rect 491986 673378 492222 673614
rect 492306 673378 492542 673614
rect 491986 673058 492222 673294
rect 492306 673058 492542 673294
rect 491986 613378 492222 613614
rect 492306 613378 492542 613614
rect 491986 613058 492222 613294
rect 492306 613058 492542 613294
rect 491986 553378 492222 553614
rect 492306 553378 492542 553614
rect 491986 553058 492222 553294
rect 492306 553058 492542 553294
rect 491986 493378 492222 493614
rect 492306 493378 492542 493614
rect 491986 493058 492222 493294
rect 492306 493058 492542 493294
rect 491986 433378 492222 433614
rect 492306 433378 492542 433614
rect 491986 433058 492222 433294
rect 492306 433058 492542 433294
rect 491986 373378 492222 373614
rect 492306 373378 492542 373614
rect 491986 373058 492222 373294
rect 492306 373058 492542 373294
rect 491986 313378 492222 313614
rect 492306 313378 492542 313614
rect 491986 313058 492222 313294
rect 492306 313058 492542 313294
rect 491986 253378 492222 253614
rect 492306 253378 492542 253614
rect 491986 253058 492222 253294
rect 492306 253058 492542 253294
rect 491986 193378 492222 193614
rect 492306 193378 492542 193614
rect 491986 193058 492222 193294
rect 492306 193058 492542 193294
rect 491986 133378 492222 133614
rect 492306 133378 492542 133614
rect 491986 133058 492222 133294
rect 492306 133058 492542 133294
rect 491986 73378 492222 73614
rect 492306 73378 492542 73614
rect 491986 73058 492222 73294
rect 492306 73058 492542 73294
rect 491986 13378 492222 13614
rect 492306 13378 492542 13614
rect 491986 13058 492222 13294
rect 492306 13058 492542 13294
rect 461986 -7302 462222 -7066
rect 462306 -7302 462542 -7066
rect 461986 -7622 462222 -7386
rect 462306 -7622 462542 -7386
rect 510826 705562 511062 705798
rect 511146 705562 511382 705798
rect 510826 705242 511062 705478
rect 511146 705242 511382 705478
rect 510826 692218 511062 692454
rect 511146 692218 511382 692454
rect 510826 691898 511062 692134
rect 511146 691898 511382 692134
rect 510826 632218 511062 632454
rect 511146 632218 511382 632454
rect 510826 631898 511062 632134
rect 511146 631898 511382 632134
rect 510826 572218 511062 572454
rect 511146 572218 511382 572454
rect 510826 571898 511062 572134
rect 511146 571898 511382 572134
rect 510826 512218 511062 512454
rect 511146 512218 511382 512454
rect 510826 511898 511062 512134
rect 511146 511898 511382 512134
rect 510826 452218 511062 452454
rect 511146 452218 511382 452454
rect 510826 451898 511062 452134
rect 511146 451898 511382 452134
rect 510826 392218 511062 392454
rect 511146 392218 511382 392454
rect 510826 391898 511062 392134
rect 511146 391898 511382 392134
rect 510826 332218 511062 332454
rect 511146 332218 511382 332454
rect 510826 331898 511062 332134
rect 511146 331898 511382 332134
rect 510826 272218 511062 272454
rect 511146 272218 511382 272454
rect 510826 271898 511062 272134
rect 511146 271898 511382 272134
rect 510826 212218 511062 212454
rect 511146 212218 511382 212454
rect 510826 211898 511062 212134
rect 511146 211898 511382 212134
rect 510826 152218 511062 152454
rect 511146 152218 511382 152454
rect 510826 151898 511062 152134
rect 511146 151898 511382 152134
rect 510826 92218 511062 92454
rect 511146 92218 511382 92454
rect 510826 91898 511062 92134
rect 511146 91898 511382 92134
rect 510826 32218 511062 32454
rect 511146 32218 511382 32454
rect 510826 31898 511062 32134
rect 511146 31898 511382 32134
rect 510826 -1542 511062 -1306
rect 511146 -1542 511382 -1306
rect 510826 -1862 511062 -1626
rect 511146 -1862 511382 -1626
rect 514546 695938 514782 696174
rect 514866 695938 515102 696174
rect 514546 695618 514782 695854
rect 514866 695618 515102 695854
rect 514546 635938 514782 636174
rect 514866 635938 515102 636174
rect 514546 635618 514782 635854
rect 514866 635618 515102 635854
rect 514546 575938 514782 576174
rect 514866 575938 515102 576174
rect 514546 575618 514782 575854
rect 514866 575618 515102 575854
rect 514546 515938 514782 516174
rect 514866 515938 515102 516174
rect 514546 515618 514782 515854
rect 514866 515618 515102 515854
rect 514546 455938 514782 456174
rect 514866 455938 515102 456174
rect 514546 455618 514782 455854
rect 514866 455618 515102 455854
rect 514546 395938 514782 396174
rect 514866 395938 515102 396174
rect 514546 395618 514782 395854
rect 514866 395618 515102 395854
rect 514546 335938 514782 336174
rect 514866 335938 515102 336174
rect 514546 335618 514782 335854
rect 514866 335618 515102 335854
rect 514546 275938 514782 276174
rect 514866 275938 515102 276174
rect 514546 275618 514782 275854
rect 514866 275618 515102 275854
rect 514546 215938 514782 216174
rect 514866 215938 515102 216174
rect 514546 215618 514782 215854
rect 514866 215618 515102 215854
rect 514546 155938 514782 156174
rect 514866 155938 515102 156174
rect 514546 155618 514782 155854
rect 514866 155618 515102 155854
rect 514546 95938 514782 96174
rect 514866 95938 515102 96174
rect 514546 95618 514782 95854
rect 514866 95618 515102 95854
rect 514546 35938 514782 36174
rect 514866 35938 515102 36174
rect 514546 35618 514782 35854
rect 514866 35618 515102 35854
rect 514546 -3462 514782 -3226
rect 514866 -3462 515102 -3226
rect 514546 -3782 514782 -3546
rect 514866 -3782 515102 -3546
rect 518266 699658 518502 699894
rect 518586 699658 518822 699894
rect 518266 699338 518502 699574
rect 518586 699338 518822 699574
rect 518266 639658 518502 639894
rect 518586 639658 518822 639894
rect 518266 639338 518502 639574
rect 518586 639338 518822 639574
rect 518266 579658 518502 579894
rect 518586 579658 518822 579894
rect 518266 579338 518502 579574
rect 518586 579338 518822 579574
rect 518266 519658 518502 519894
rect 518586 519658 518822 519894
rect 518266 519338 518502 519574
rect 518586 519338 518822 519574
rect 518266 459658 518502 459894
rect 518586 459658 518822 459894
rect 518266 459338 518502 459574
rect 518586 459338 518822 459574
rect 518266 399658 518502 399894
rect 518586 399658 518822 399894
rect 518266 399338 518502 399574
rect 518586 399338 518822 399574
rect 518266 339658 518502 339894
rect 518586 339658 518822 339894
rect 518266 339338 518502 339574
rect 518586 339338 518822 339574
rect 518266 279658 518502 279894
rect 518586 279658 518822 279894
rect 518266 279338 518502 279574
rect 518586 279338 518822 279574
rect 518266 219658 518502 219894
rect 518586 219658 518822 219894
rect 518266 219338 518502 219574
rect 518586 219338 518822 219574
rect 518266 159658 518502 159894
rect 518586 159658 518822 159894
rect 518266 159338 518502 159574
rect 518586 159338 518822 159574
rect 518266 99658 518502 99894
rect 518586 99658 518822 99894
rect 518266 99338 518502 99574
rect 518586 99338 518822 99574
rect 518266 39658 518502 39894
rect 518586 39658 518822 39894
rect 518266 39338 518502 39574
rect 518586 39338 518822 39574
rect 518266 -5382 518502 -5146
rect 518586 -5382 518822 -5146
rect 518266 -5702 518502 -5466
rect 518586 -5702 518822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 551986 710362 552222 710598
rect 552306 710362 552542 710598
rect 551986 710042 552222 710278
rect 552306 710042 552542 710278
rect 548266 708442 548502 708678
rect 548586 708442 548822 708678
rect 548266 708122 548502 708358
rect 548586 708122 548822 708358
rect 544546 706522 544782 706758
rect 544866 706522 545102 706758
rect 544546 706202 544782 706438
rect 544866 706202 545102 706438
rect 521986 643378 522222 643614
rect 522306 643378 522542 643614
rect 521986 643058 522222 643294
rect 522306 643058 522542 643294
rect 521986 583378 522222 583614
rect 522306 583378 522542 583614
rect 521986 583058 522222 583294
rect 522306 583058 522542 583294
rect 521986 523378 522222 523614
rect 522306 523378 522542 523614
rect 521986 523058 522222 523294
rect 522306 523058 522542 523294
rect 521986 463378 522222 463614
rect 522306 463378 522542 463614
rect 521986 463058 522222 463294
rect 522306 463058 522542 463294
rect 521986 403378 522222 403614
rect 522306 403378 522542 403614
rect 521986 403058 522222 403294
rect 522306 403058 522542 403294
rect 521986 343378 522222 343614
rect 522306 343378 522542 343614
rect 521986 343058 522222 343294
rect 522306 343058 522542 343294
rect 521986 283378 522222 283614
rect 522306 283378 522542 283614
rect 521986 283058 522222 283294
rect 522306 283058 522542 283294
rect 521986 223378 522222 223614
rect 522306 223378 522542 223614
rect 521986 223058 522222 223294
rect 522306 223058 522542 223294
rect 521986 163378 522222 163614
rect 522306 163378 522542 163614
rect 521986 163058 522222 163294
rect 522306 163058 522542 163294
rect 521986 103378 522222 103614
rect 522306 103378 522542 103614
rect 521986 103058 522222 103294
rect 522306 103058 522542 103294
rect 521986 43378 522222 43614
rect 522306 43378 522542 43614
rect 521986 43058 522222 43294
rect 522306 43058 522542 43294
rect 491986 -6342 492222 -6106
rect 492306 -6342 492542 -6106
rect 491986 -6662 492222 -6426
rect 492306 -6662 492542 -6426
rect 540826 704602 541062 704838
rect 541146 704602 541382 704838
rect 540826 704282 541062 704518
rect 541146 704282 541382 704518
rect 540826 662218 541062 662454
rect 541146 662218 541382 662454
rect 540826 661898 541062 662134
rect 541146 661898 541382 662134
rect 540826 602218 541062 602454
rect 541146 602218 541382 602454
rect 540826 601898 541062 602134
rect 541146 601898 541382 602134
rect 540826 542218 541062 542454
rect 541146 542218 541382 542454
rect 540826 541898 541062 542134
rect 541146 541898 541382 542134
rect 540826 482218 541062 482454
rect 541146 482218 541382 482454
rect 540826 481898 541062 482134
rect 541146 481898 541382 482134
rect 540826 422218 541062 422454
rect 541146 422218 541382 422454
rect 540826 421898 541062 422134
rect 541146 421898 541382 422134
rect 540826 362218 541062 362454
rect 541146 362218 541382 362454
rect 540826 361898 541062 362134
rect 541146 361898 541382 362134
rect 540826 302218 541062 302454
rect 541146 302218 541382 302454
rect 540826 301898 541062 302134
rect 541146 301898 541382 302134
rect 540826 242218 541062 242454
rect 541146 242218 541382 242454
rect 540826 241898 541062 242134
rect 541146 241898 541382 242134
rect 540826 182218 541062 182454
rect 541146 182218 541382 182454
rect 540826 181898 541062 182134
rect 541146 181898 541382 182134
rect 540826 122218 541062 122454
rect 541146 122218 541382 122454
rect 540826 121898 541062 122134
rect 541146 121898 541382 122134
rect 540826 62218 541062 62454
rect 541146 62218 541382 62454
rect 540826 61898 541062 62134
rect 541146 61898 541382 62134
rect 540826 2218 541062 2454
rect 541146 2218 541382 2454
rect 540826 1898 541062 2134
rect 541146 1898 541382 2134
rect 540826 -582 541062 -346
rect 541146 -582 541382 -346
rect 540826 -902 541062 -666
rect 541146 -902 541382 -666
rect 544546 665938 544782 666174
rect 544866 665938 545102 666174
rect 544546 665618 544782 665854
rect 544866 665618 545102 665854
rect 544546 605938 544782 606174
rect 544866 605938 545102 606174
rect 544546 605618 544782 605854
rect 544866 605618 545102 605854
rect 544546 545938 544782 546174
rect 544866 545938 545102 546174
rect 544546 545618 544782 545854
rect 544866 545618 545102 545854
rect 544546 485938 544782 486174
rect 544866 485938 545102 486174
rect 544546 485618 544782 485854
rect 544866 485618 545102 485854
rect 544546 425938 544782 426174
rect 544866 425938 545102 426174
rect 544546 425618 544782 425854
rect 544866 425618 545102 425854
rect 544546 365938 544782 366174
rect 544866 365938 545102 366174
rect 544546 365618 544782 365854
rect 544866 365618 545102 365854
rect 544546 305938 544782 306174
rect 544866 305938 545102 306174
rect 544546 305618 544782 305854
rect 544866 305618 545102 305854
rect 544546 245938 544782 246174
rect 544866 245938 545102 246174
rect 544546 245618 544782 245854
rect 544866 245618 545102 245854
rect 544546 185938 544782 186174
rect 544866 185938 545102 186174
rect 544546 185618 544782 185854
rect 544866 185618 545102 185854
rect 544546 125938 544782 126174
rect 544866 125938 545102 126174
rect 544546 125618 544782 125854
rect 544866 125618 545102 125854
rect 544546 65938 544782 66174
rect 544866 65938 545102 66174
rect 544546 65618 544782 65854
rect 544866 65618 545102 65854
rect 544546 5938 544782 6174
rect 544866 5938 545102 6174
rect 544546 5618 544782 5854
rect 544866 5618 545102 5854
rect 544546 -2502 544782 -2266
rect 544866 -2502 545102 -2266
rect 544546 -2822 544782 -2586
rect 544866 -2822 545102 -2586
rect 548266 669658 548502 669894
rect 548586 669658 548822 669894
rect 548266 669338 548502 669574
rect 548586 669338 548822 669574
rect 548266 609658 548502 609894
rect 548586 609658 548822 609894
rect 548266 609338 548502 609574
rect 548586 609338 548822 609574
rect 548266 549658 548502 549894
rect 548586 549658 548822 549894
rect 548266 549338 548502 549574
rect 548586 549338 548822 549574
rect 548266 489658 548502 489894
rect 548586 489658 548822 489894
rect 548266 489338 548502 489574
rect 548586 489338 548822 489574
rect 548266 429658 548502 429894
rect 548586 429658 548822 429894
rect 548266 429338 548502 429574
rect 548586 429338 548822 429574
rect 548266 369658 548502 369894
rect 548586 369658 548822 369894
rect 548266 369338 548502 369574
rect 548586 369338 548822 369574
rect 548266 309658 548502 309894
rect 548586 309658 548822 309894
rect 548266 309338 548502 309574
rect 548586 309338 548822 309574
rect 548266 249658 548502 249894
rect 548586 249658 548822 249894
rect 548266 249338 548502 249574
rect 548586 249338 548822 249574
rect 548266 189658 548502 189894
rect 548586 189658 548822 189894
rect 548266 189338 548502 189574
rect 548586 189338 548822 189574
rect 548266 129658 548502 129894
rect 548586 129658 548822 129894
rect 548266 129338 548502 129574
rect 548586 129338 548822 129574
rect 548266 69658 548502 69894
rect 548586 69658 548822 69894
rect 548266 69338 548502 69574
rect 548586 69338 548822 69574
rect 548266 9658 548502 9894
rect 548586 9658 548822 9894
rect 548266 9338 548502 9574
rect 548586 9338 548822 9574
rect 548266 -4422 548502 -4186
rect 548586 -4422 548822 -4186
rect 548266 -4742 548502 -4506
rect 548586 -4742 548822 -4506
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 578266 709402 578502 709638
rect 578586 709402 578822 709638
rect 578266 709082 578502 709318
rect 578586 709082 578822 709318
rect 574546 707482 574782 707718
rect 574866 707482 575102 707718
rect 574546 707162 574782 707398
rect 574866 707162 575102 707398
rect 551986 673378 552222 673614
rect 552306 673378 552542 673614
rect 551986 673058 552222 673294
rect 552306 673058 552542 673294
rect 551986 613378 552222 613614
rect 552306 613378 552542 613614
rect 551986 613058 552222 613294
rect 552306 613058 552542 613294
rect 551986 553378 552222 553614
rect 552306 553378 552542 553614
rect 551986 553058 552222 553294
rect 552306 553058 552542 553294
rect 551986 493378 552222 493614
rect 552306 493378 552542 493614
rect 551986 493058 552222 493294
rect 552306 493058 552542 493294
rect 551986 433378 552222 433614
rect 552306 433378 552542 433614
rect 551986 433058 552222 433294
rect 552306 433058 552542 433294
rect 551986 373378 552222 373614
rect 552306 373378 552542 373614
rect 551986 373058 552222 373294
rect 552306 373058 552542 373294
rect 551986 313378 552222 313614
rect 552306 313378 552542 313614
rect 551986 313058 552222 313294
rect 552306 313058 552542 313294
rect 551986 253378 552222 253614
rect 552306 253378 552542 253614
rect 551986 253058 552222 253294
rect 552306 253058 552542 253294
rect 551986 193378 552222 193614
rect 552306 193378 552542 193614
rect 551986 193058 552222 193294
rect 552306 193058 552542 193294
rect 551986 133378 552222 133614
rect 552306 133378 552542 133614
rect 551986 133058 552222 133294
rect 552306 133058 552542 133294
rect 551986 73378 552222 73614
rect 552306 73378 552542 73614
rect 551986 73058 552222 73294
rect 552306 73058 552542 73294
rect 551986 13378 552222 13614
rect 552306 13378 552542 13614
rect 551986 13058 552222 13294
rect 552306 13058 552542 13294
rect 521986 -7302 522222 -7066
rect 522306 -7302 522542 -7066
rect 521986 -7622 522222 -7386
rect 522306 -7622 522542 -7386
rect 570826 705562 571062 705798
rect 571146 705562 571382 705798
rect 570826 705242 571062 705478
rect 571146 705242 571382 705478
rect 570826 692218 571062 692454
rect 571146 692218 571382 692454
rect 570826 691898 571062 692134
rect 571146 691898 571382 692134
rect 570826 632218 571062 632454
rect 571146 632218 571382 632454
rect 570826 631898 571062 632134
rect 571146 631898 571382 632134
rect 570826 572218 571062 572454
rect 571146 572218 571382 572454
rect 570826 571898 571062 572134
rect 571146 571898 571382 572134
rect 570826 512218 571062 512454
rect 571146 512218 571382 512454
rect 570826 511898 571062 512134
rect 571146 511898 571382 512134
rect 570826 452218 571062 452454
rect 571146 452218 571382 452454
rect 570826 451898 571062 452134
rect 571146 451898 571382 452134
rect 570826 392218 571062 392454
rect 571146 392218 571382 392454
rect 570826 391898 571062 392134
rect 571146 391898 571382 392134
rect 570826 332218 571062 332454
rect 571146 332218 571382 332454
rect 570826 331898 571062 332134
rect 571146 331898 571382 332134
rect 570826 272218 571062 272454
rect 571146 272218 571382 272454
rect 570826 271898 571062 272134
rect 571146 271898 571382 272134
rect 570826 212218 571062 212454
rect 571146 212218 571382 212454
rect 570826 211898 571062 212134
rect 571146 211898 571382 212134
rect 570826 152218 571062 152454
rect 571146 152218 571382 152454
rect 570826 151898 571062 152134
rect 571146 151898 571382 152134
rect 570826 92218 571062 92454
rect 571146 92218 571382 92454
rect 570826 91898 571062 92134
rect 571146 91898 571382 92134
rect 570826 32218 571062 32454
rect 571146 32218 571382 32454
rect 570826 31898 571062 32134
rect 571146 31898 571382 32134
rect 570826 -1542 571062 -1306
rect 571146 -1542 571382 -1306
rect 570826 -1862 571062 -1626
rect 571146 -1862 571382 -1626
rect 574546 695938 574782 696174
rect 574866 695938 575102 696174
rect 574546 695618 574782 695854
rect 574866 695618 575102 695854
rect 574546 635938 574782 636174
rect 574866 635938 575102 636174
rect 574546 635618 574782 635854
rect 574866 635618 575102 635854
rect 574546 575938 574782 576174
rect 574866 575938 575102 576174
rect 574546 575618 574782 575854
rect 574866 575618 575102 575854
rect 574546 515938 574782 516174
rect 574866 515938 575102 516174
rect 574546 515618 574782 515854
rect 574866 515618 575102 515854
rect 574546 455938 574782 456174
rect 574866 455938 575102 456174
rect 574546 455618 574782 455854
rect 574866 455618 575102 455854
rect 574546 395938 574782 396174
rect 574866 395938 575102 396174
rect 574546 395618 574782 395854
rect 574866 395618 575102 395854
rect 574546 335938 574782 336174
rect 574866 335938 575102 336174
rect 574546 335618 574782 335854
rect 574866 335618 575102 335854
rect 574546 275938 574782 276174
rect 574866 275938 575102 276174
rect 574546 275618 574782 275854
rect 574866 275618 575102 275854
rect 574546 215938 574782 216174
rect 574866 215938 575102 216174
rect 574546 215618 574782 215854
rect 574866 215618 575102 215854
rect 574546 155938 574782 156174
rect 574866 155938 575102 156174
rect 574546 155618 574782 155854
rect 574866 155618 575102 155854
rect 574546 95938 574782 96174
rect 574866 95938 575102 96174
rect 574546 95618 574782 95854
rect 574866 95618 575102 95854
rect 574546 35938 574782 36174
rect 574866 35938 575102 36174
rect 574546 35618 574782 35854
rect 574866 35618 575102 35854
rect 574546 -3462 574782 -3226
rect 574866 -3462 575102 -3226
rect 574546 -3782 574782 -3546
rect 574866 -3782 575102 -3546
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 578266 699658 578502 699894
rect 578586 699658 578822 699894
rect 578266 699338 578502 699574
rect 578586 699338 578822 699574
rect 578266 639658 578502 639894
rect 578586 639658 578822 639894
rect 578266 639338 578502 639574
rect 578586 639338 578822 639574
rect 578266 579658 578502 579894
rect 578586 579658 578822 579894
rect 578266 579338 578502 579574
rect 578586 579338 578822 579574
rect 578266 519658 578502 519894
rect 578586 519658 578822 519894
rect 578266 519338 578502 519574
rect 578586 519338 578822 519574
rect 578266 459658 578502 459894
rect 578586 459658 578822 459894
rect 578266 459338 578502 459574
rect 578586 459338 578822 459574
rect 578266 399658 578502 399894
rect 578586 399658 578822 399894
rect 578266 399338 578502 399574
rect 578586 399338 578822 399574
rect 578266 339658 578502 339894
rect 578586 339658 578822 339894
rect 578266 339338 578502 339574
rect 578586 339338 578822 339574
rect 578266 279658 578502 279894
rect 578586 279658 578822 279894
rect 578266 279338 578502 279574
rect 578586 279338 578822 279574
rect 578266 219658 578502 219894
rect 578586 219658 578822 219894
rect 578266 219338 578502 219574
rect 578586 219338 578822 219574
rect 578266 159658 578502 159894
rect 578586 159658 578822 159894
rect 578266 159338 578502 159574
rect 578586 159338 578822 159574
rect 578266 99658 578502 99894
rect 578586 99658 578822 99894
rect 578266 99338 578502 99574
rect 578586 99338 578822 99574
rect 578266 39658 578502 39894
rect 578586 39658 578822 39894
rect 578266 39338 578502 39574
rect 578586 39338 578822 39574
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 662218 585578 662454
rect 585662 662218 585898 662454
rect 585342 661898 585578 662134
rect 585662 661898 585898 662134
rect 585342 602218 585578 602454
rect 585662 602218 585898 602454
rect 585342 601898 585578 602134
rect 585662 601898 585898 602134
rect 585342 542218 585578 542454
rect 585662 542218 585898 542454
rect 585342 541898 585578 542134
rect 585662 541898 585898 542134
rect 585342 482218 585578 482454
rect 585662 482218 585898 482454
rect 585342 481898 585578 482134
rect 585662 481898 585898 482134
rect 585342 422218 585578 422454
rect 585662 422218 585898 422454
rect 585342 421898 585578 422134
rect 585662 421898 585898 422134
rect 585342 362218 585578 362454
rect 585662 362218 585898 362454
rect 585342 361898 585578 362134
rect 585662 361898 585898 362134
rect 585342 302218 585578 302454
rect 585662 302218 585898 302454
rect 585342 301898 585578 302134
rect 585662 301898 585898 302134
rect 585342 242218 585578 242454
rect 585662 242218 585898 242454
rect 585342 241898 585578 242134
rect 585662 241898 585898 242134
rect 585342 182218 585578 182454
rect 585662 182218 585898 182454
rect 585342 181898 585578 182134
rect 585662 181898 585898 182134
rect 585342 122218 585578 122454
rect 585662 122218 585898 122454
rect 585342 121898 585578 122134
rect 585662 121898 585898 122134
rect 585342 62218 585578 62454
rect 585662 62218 585898 62454
rect 585342 61898 585578 62134
rect 585662 61898 585898 62134
rect 585342 2218 585578 2454
rect 585662 2218 585898 2454
rect 585342 1898 585578 2134
rect 585662 1898 585898 2134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 692218 586538 692454
rect 586622 692218 586858 692454
rect 586302 691898 586538 692134
rect 586622 691898 586858 692134
rect 586302 632218 586538 632454
rect 586622 632218 586858 632454
rect 586302 631898 586538 632134
rect 586622 631898 586858 632134
rect 586302 572218 586538 572454
rect 586622 572218 586858 572454
rect 586302 571898 586538 572134
rect 586622 571898 586858 572134
rect 586302 512218 586538 512454
rect 586622 512218 586858 512454
rect 586302 511898 586538 512134
rect 586622 511898 586858 512134
rect 586302 452218 586538 452454
rect 586622 452218 586858 452454
rect 586302 451898 586538 452134
rect 586622 451898 586858 452134
rect 586302 392218 586538 392454
rect 586622 392218 586858 392454
rect 586302 391898 586538 392134
rect 586622 391898 586858 392134
rect 586302 332218 586538 332454
rect 586622 332218 586858 332454
rect 586302 331898 586538 332134
rect 586622 331898 586858 332134
rect 586302 272218 586538 272454
rect 586622 272218 586858 272454
rect 586302 271898 586538 272134
rect 586622 271898 586858 272134
rect 586302 212218 586538 212454
rect 586622 212218 586858 212454
rect 586302 211898 586538 212134
rect 586622 211898 586858 212134
rect 586302 152218 586538 152454
rect 586622 152218 586858 152454
rect 586302 151898 586538 152134
rect 586622 151898 586858 152134
rect 586302 92218 586538 92454
rect 586622 92218 586858 92454
rect 586302 91898 586538 92134
rect 586622 91898 586858 92134
rect 586302 32218 586538 32454
rect 586622 32218 586858 32454
rect 586302 31898 586538 32134
rect 586622 31898 586858 32134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 665938 587498 666174
rect 587582 665938 587818 666174
rect 587262 665618 587498 665854
rect 587582 665618 587818 665854
rect 587262 605938 587498 606174
rect 587582 605938 587818 606174
rect 587262 605618 587498 605854
rect 587582 605618 587818 605854
rect 587262 545938 587498 546174
rect 587582 545938 587818 546174
rect 587262 545618 587498 545854
rect 587582 545618 587818 545854
rect 587262 485938 587498 486174
rect 587582 485938 587818 486174
rect 587262 485618 587498 485854
rect 587582 485618 587818 485854
rect 587262 425938 587498 426174
rect 587582 425938 587818 426174
rect 587262 425618 587498 425854
rect 587582 425618 587818 425854
rect 587262 365938 587498 366174
rect 587582 365938 587818 366174
rect 587262 365618 587498 365854
rect 587582 365618 587818 365854
rect 587262 305938 587498 306174
rect 587582 305938 587818 306174
rect 587262 305618 587498 305854
rect 587582 305618 587818 305854
rect 587262 245938 587498 246174
rect 587582 245938 587818 246174
rect 587262 245618 587498 245854
rect 587582 245618 587818 245854
rect 587262 185938 587498 186174
rect 587582 185938 587818 186174
rect 587262 185618 587498 185854
rect 587582 185618 587818 185854
rect 587262 125938 587498 126174
rect 587582 125938 587818 126174
rect 587262 125618 587498 125854
rect 587582 125618 587818 125854
rect 587262 65938 587498 66174
rect 587582 65938 587818 66174
rect 587262 65618 587498 65854
rect 587582 65618 587818 65854
rect 587262 5938 587498 6174
rect 587582 5938 587818 6174
rect 587262 5618 587498 5854
rect 587582 5618 587818 5854
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 695938 588458 696174
rect 588542 695938 588778 696174
rect 588222 695618 588458 695854
rect 588542 695618 588778 695854
rect 588222 635938 588458 636174
rect 588542 635938 588778 636174
rect 588222 635618 588458 635854
rect 588542 635618 588778 635854
rect 588222 575938 588458 576174
rect 588542 575938 588778 576174
rect 588222 575618 588458 575854
rect 588542 575618 588778 575854
rect 588222 515938 588458 516174
rect 588542 515938 588778 516174
rect 588222 515618 588458 515854
rect 588542 515618 588778 515854
rect 588222 455938 588458 456174
rect 588542 455938 588778 456174
rect 588222 455618 588458 455854
rect 588542 455618 588778 455854
rect 588222 395938 588458 396174
rect 588542 395938 588778 396174
rect 588222 395618 588458 395854
rect 588542 395618 588778 395854
rect 588222 335938 588458 336174
rect 588542 335938 588778 336174
rect 588222 335618 588458 335854
rect 588542 335618 588778 335854
rect 588222 275938 588458 276174
rect 588542 275938 588778 276174
rect 588222 275618 588458 275854
rect 588542 275618 588778 275854
rect 588222 215938 588458 216174
rect 588542 215938 588778 216174
rect 588222 215618 588458 215854
rect 588542 215618 588778 215854
rect 588222 155938 588458 156174
rect 588542 155938 588778 156174
rect 588222 155618 588458 155854
rect 588542 155618 588778 155854
rect 588222 95938 588458 96174
rect 588542 95938 588778 96174
rect 588222 95618 588458 95854
rect 588542 95618 588778 95854
rect 588222 35938 588458 36174
rect 588542 35938 588778 36174
rect 588222 35618 588458 35854
rect 588542 35618 588778 35854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669658 589418 669894
rect 589502 669658 589738 669894
rect 589182 669338 589418 669574
rect 589502 669338 589738 669574
rect 589182 609658 589418 609894
rect 589502 609658 589738 609894
rect 589182 609338 589418 609574
rect 589502 609338 589738 609574
rect 589182 549658 589418 549894
rect 589502 549658 589738 549894
rect 589182 549338 589418 549574
rect 589502 549338 589738 549574
rect 589182 489658 589418 489894
rect 589502 489658 589738 489894
rect 589182 489338 589418 489574
rect 589502 489338 589738 489574
rect 589182 429658 589418 429894
rect 589502 429658 589738 429894
rect 589182 429338 589418 429574
rect 589502 429338 589738 429574
rect 589182 369658 589418 369894
rect 589502 369658 589738 369894
rect 589182 369338 589418 369574
rect 589502 369338 589738 369574
rect 589182 309658 589418 309894
rect 589502 309658 589738 309894
rect 589182 309338 589418 309574
rect 589502 309338 589738 309574
rect 589182 249658 589418 249894
rect 589502 249658 589738 249894
rect 589182 249338 589418 249574
rect 589502 249338 589738 249574
rect 589182 189658 589418 189894
rect 589502 189658 589738 189894
rect 589182 189338 589418 189574
rect 589502 189338 589738 189574
rect 589182 129658 589418 129894
rect 589502 129658 589738 129894
rect 589182 129338 589418 129574
rect 589502 129338 589738 129574
rect 589182 69658 589418 69894
rect 589502 69658 589738 69894
rect 589182 69338 589418 69574
rect 589502 69338 589738 69574
rect 589182 9658 589418 9894
rect 589502 9658 589738 9894
rect 589182 9338 589418 9574
rect 589502 9338 589738 9574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 699658 590378 699894
rect 590462 699658 590698 699894
rect 590142 699338 590378 699574
rect 590462 699338 590698 699574
rect 590142 639658 590378 639894
rect 590462 639658 590698 639894
rect 590142 639338 590378 639574
rect 590462 639338 590698 639574
rect 590142 579658 590378 579894
rect 590462 579658 590698 579894
rect 590142 579338 590378 579574
rect 590462 579338 590698 579574
rect 590142 519658 590378 519894
rect 590462 519658 590698 519894
rect 590142 519338 590378 519574
rect 590462 519338 590698 519574
rect 590142 459658 590378 459894
rect 590462 459658 590698 459894
rect 590142 459338 590378 459574
rect 590462 459338 590698 459574
rect 590142 399658 590378 399894
rect 590462 399658 590698 399894
rect 590142 399338 590378 399574
rect 590462 399338 590698 399574
rect 590142 339658 590378 339894
rect 590462 339658 590698 339894
rect 590142 339338 590378 339574
rect 590462 339338 590698 339574
rect 590142 279658 590378 279894
rect 590462 279658 590698 279894
rect 590142 279338 590378 279574
rect 590462 279338 590698 279574
rect 590142 219658 590378 219894
rect 590462 219658 590698 219894
rect 590142 219338 590378 219574
rect 590462 219338 590698 219574
rect 590142 159658 590378 159894
rect 590462 159658 590698 159894
rect 590142 159338 590378 159574
rect 590462 159338 590698 159574
rect 590142 99658 590378 99894
rect 590462 99658 590698 99894
rect 590142 99338 590378 99574
rect 590462 99338 590698 99574
rect 590142 39658 590378 39894
rect 590462 39658 590698 39894
rect 590142 39338 590378 39574
rect 590462 39338 590698 39574
rect 578266 -5382 578502 -5146
rect 578586 -5382 578822 -5146
rect 578266 -5702 578502 -5466
rect 578586 -5702 578822 -5466
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673378 591338 673614
rect 591422 673378 591658 673614
rect 591102 673058 591338 673294
rect 591422 673058 591658 673294
rect 591102 613378 591338 613614
rect 591422 613378 591658 613614
rect 591102 613058 591338 613294
rect 591422 613058 591658 613294
rect 591102 553378 591338 553614
rect 591422 553378 591658 553614
rect 591102 553058 591338 553294
rect 591422 553058 591658 553294
rect 591102 493378 591338 493614
rect 591422 493378 591658 493614
rect 591102 493058 591338 493294
rect 591422 493058 591658 493294
rect 591102 433378 591338 433614
rect 591422 433378 591658 433614
rect 591102 433058 591338 433294
rect 591422 433058 591658 433294
rect 591102 373378 591338 373614
rect 591422 373378 591658 373614
rect 591102 373058 591338 373294
rect 591422 373058 591658 373294
rect 591102 313378 591338 313614
rect 591422 313378 591658 313614
rect 591102 313058 591338 313294
rect 591422 313058 591658 313294
rect 591102 253378 591338 253614
rect 591422 253378 591658 253614
rect 591102 253058 591338 253294
rect 591422 253058 591658 253294
rect 591102 193378 591338 193614
rect 591422 193378 591658 193614
rect 591102 193058 591338 193294
rect 591422 193058 591658 193294
rect 591102 133378 591338 133614
rect 591422 133378 591658 133614
rect 591102 133058 591338 133294
rect 591422 133058 591658 133294
rect 591102 73378 591338 73614
rect 591422 73378 591658 73614
rect 591102 73058 591338 73294
rect 591422 73058 591658 73294
rect 591102 13378 591338 13614
rect 591422 13378 591658 13614
rect 591102 13058 591338 13294
rect 591422 13058 591658 13294
rect 551986 -6342 552222 -6106
rect 552306 -6342 552542 -6106
rect 551986 -6662 552222 -6426
rect 552306 -6662 552542 -6426
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 643378 592298 643614
rect 592382 643378 592618 643614
rect 592062 643058 592298 643294
rect 592382 643058 592618 643294
rect 592062 583378 592298 583614
rect 592382 583378 592618 583614
rect 592062 583058 592298 583294
rect 592382 583058 592618 583294
rect 592062 523378 592298 523614
rect 592382 523378 592618 523614
rect 592062 523058 592298 523294
rect 592382 523058 592618 523294
rect 592062 463378 592298 463614
rect 592382 463378 592618 463614
rect 592062 463058 592298 463294
rect 592382 463058 592618 463294
rect 592062 403378 592298 403614
rect 592382 403378 592618 403614
rect 592062 403058 592298 403294
rect 592382 403058 592618 403294
rect 592062 343378 592298 343614
rect 592382 343378 592618 343614
rect 592062 343058 592298 343294
rect 592382 343058 592618 343294
rect 592062 283378 592298 283614
rect 592382 283378 592618 283614
rect 592062 283058 592298 283294
rect 592382 283058 592618 283294
rect 592062 223378 592298 223614
rect 592382 223378 592618 223614
rect 592062 223058 592298 223294
rect 592382 223058 592618 223294
rect 592062 163378 592298 163614
rect 592382 163378 592618 163614
rect 592062 163058 592298 163294
rect 592382 163058 592618 163294
rect 592062 103378 592298 103614
rect 592382 103378 592618 103614
rect 592062 103058 592298 103294
rect 592382 103058 592618 103294
rect 592062 43378 592298 43614
rect 592382 43378 592618 43614
rect 592062 43058 592298 43294
rect 592382 43058 592618 43294
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 41986 711558
rect 42222 711322 42306 711558
rect 42542 711322 101986 711558
rect 102222 711322 102306 711558
rect 102542 711322 161986 711558
rect 162222 711322 162306 711558
rect 162542 711322 221986 711558
rect 222222 711322 222306 711558
rect 222542 711322 281986 711558
rect 282222 711322 282306 711558
rect 282542 711322 341986 711558
rect 342222 711322 342306 711558
rect 342542 711322 401986 711558
rect 402222 711322 402306 711558
rect 402542 711322 461986 711558
rect 462222 711322 462306 711558
rect 462542 711322 521986 711558
rect 522222 711322 522306 711558
rect 522542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 41986 711238
rect 42222 711002 42306 711238
rect 42542 711002 101986 711238
rect 102222 711002 102306 711238
rect 102542 711002 161986 711238
rect 162222 711002 162306 711238
rect 162542 711002 221986 711238
rect 222222 711002 222306 711238
rect 222542 711002 281986 711238
rect 282222 711002 282306 711238
rect 282542 711002 341986 711238
rect 342222 711002 342306 711238
rect 342542 711002 401986 711238
rect 402222 711002 402306 711238
rect 402542 711002 461986 711238
rect 462222 711002 462306 711238
rect 462542 711002 521986 711238
rect 522222 711002 522306 711238
rect 522542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 11986 710598
rect 12222 710362 12306 710598
rect 12542 710362 71986 710598
rect 72222 710362 72306 710598
rect 72542 710362 131986 710598
rect 132222 710362 132306 710598
rect 132542 710362 191986 710598
rect 192222 710362 192306 710598
rect 192542 710362 251986 710598
rect 252222 710362 252306 710598
rect 252542 710362 311986 710598
rect 312222 710362 312306 710598
rect 312542 710362 371986 710598
rect 372222 710362 372306 710598
rect 372542 710362 431986 710598
rect 432222 710362 432306 710598
rect 432542 710362 491986 710598
rect 492222 710362 492306 710598
rect 492542 710362 551986 710598
rect 552222 710362 552306 710598
rect 552542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 11986 710278
rect 12222 710042 12306 710278
rect 12542 710042 71986 710278
rect 72222 710042 72306 710278
rect 72542 710042 131986 710278
rect 132222 710042 132306 710278
rect 132542 710042 191986 710278
rect 192222 710042 192306 710278
rect 192542 710042 251986 710278
rect 252222 710042 252306 710278
rect 252542 710042 311986 710278
rect 312222 710042 312306 710278
rect 312542 710042 371986 710278
rect 372222 710042 372306 710278
rect 372542 710042 431986 710278
rect 432222 710042 432306 710278
rect 432542 710042 491986 710278
rect 492222 710042 492306 710278
rect 492542 710042 551986 710278
rect 552222 710042 552306 710278
rect 552542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 38266 709638
rect 38502 709402 38586 709638
rect 38822 709402 98266 709638
rect 98502 709402 98586 709638
rect 98822 709402 158266 709638
rect 158502 709402 158586 709638
rect 158822 709402 218266 709638
rect 218502 709402 218586 709638
rect 218822 709402 278266 709638
rect 278502 709402 278586 709638
rect 278822 709402 338266 709638
rect 338502 709402 338586 709638
rect 338822 709402 398266 709638
rect 398502 709402 398586 709638
rect 398822 709402 458266 709638
rect 458502 709402 458586 709638
rect 458822 709402 518266 709638
rect 518502 709402 518586 709638
rect 518822 709402 578266 709638
rect 578502 709402 578586 709638
rect 578822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 38266 709318
rect 38502 709082 38586 709318
rect 38822 709082 98266 709318
rect 98502 709082 98586 709318
rect 98822 709082 158266 709318
rect 158502 709082 158586 709318
rect 158822 709082 218266 709318
rect 218502 709082 218586 709318
rect 218822 709082 278266 709318
rect 278502 709082 278586 709318
rect 278822 709082 338266 709318
rect 338502 709082 338586 709318
rect 338822 709082 398266 709318
rect 398502 709082 398586 709318
rect 398822 709082 458266 709318
rect 458502 709082 458586 709318
rect 458822 709082 518266 709318
rect 518502 709082 518586 709318
rect 518822 709082 578266 709318
rect 578502 709082 578586 709318
rect 578822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 8266 708678
rect 8502 708442 8586 708678
rect 8822 708442 68266 708678
rect 68502 708442 68586 708678
rect 68822 708442 128266 708678
rect 128502 708442 128586 708678
rect 128822 708442 188266 708678
rect 188502 708442 188586 708678
rect 188822 708442 248266 708678
rect 248502 708442 248586 708678
rect 248822 708442 308266 708678
rect 308502 708442 308586 708678
rect 308822 708442 368266 708678
rect 368502 708442 368586 708678
rect 368822 708442 428266 708678
rect 428502 708442 428586 708678
rect 428822 708442 488266 708678
rect 488502 708442 488586 708678
rect 488822 708442 548266 708678
rect 548502 708442 548586 708678
rect 548822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 8266 708358
rect 8502 708122 8586 708358
rect 8822 708122 68266 708358
rect 68502 708122 68586 708358
rect 68822 708122 128266 708358
rect 128502 708122 128586 708358
rect 128822 708122 188266 708358
rect 188502 708122 188586 708358
rect 188822 708122 248266 708358
rect 248502 708122 248586 708358
rect 248822 708122 308266 708358
rect 308502 708122 308586 708358
rect 308822 708122 368266 708358
rect 368502 708122 368586 708358
rect 368822 708122 428266 708358
rect 428502 708122 428586 708358
rect 428822 708122 488266 708358
rect 488502 708122 488586 708358
rect 488822 708122 548266 708358
rect 548502 708122 548586 708358
rect 548822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 34546 707718
rect 34782 707482 34866 707718
rect 35102 707482 94546 707718
rect 94782 707482 94866 707718
rect 95102 707482 154546 707718
rect 154782 707482 154866 707718
rect 155102 707482 214546 707718
rect 214782 707482 214866 707718
rect 215102 707482 274546 707718
rect 274782 707482 274866 707718
rect 275102 707482 334546 707718
rect 334782 707482 334866 707718
rect 335102 707482 394546 707718
rect 394782 707482 394866 707718
rect 395102 707482 454546 707718
rect 454782 707482 454866 707718
rect 455102 707482 514546 707718
rect 514782 707482 514866 707718
rect 515102 707482 574546 707718
rect 574782 707482 574866 707718
rect 575102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 34546 707398
rect 34782 707162 34866 707398
rect 35102 707162 94546 707398
rect 94782 707162 94866 707398
rect 95102 707162 154546 707398
rect 154782 707162 154866 707398
rect 155102 707162 214546 707398
rect 214782 707162 214866 707398
rect 215102 707162 274546 707398
rect 274782 707162 274866 707398
rect 275102 707162 334546 707398
rect 334782 707162 334866 707398
rect 335102 707162 394546 707398
rect 394782 707162 394866 707398
rect 395102 707162 454546 707398
rect 454782 707162 454866 707398
rect 455102 707162 514546 707398
rect 514782 707162 514866 707398
rect 515102 707162 574546 707398
rect 574782 707162 574866 707398
rect 575102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 4546 706758
rect 4782 706522 4866 706758
rect 5102 706522 64546 706758
rect 64782 706522 64866 706758
rect 65102 706522 124546 706758
rect 124782 706522 124866 706758
rect 125102 706522 184546 706758
rect 184782 706522 184866 706758
rect 185102 706522 244546 706758
rect 244782 706522 244866 706758
rect 245102 706522 304546 706758
rect 304782 706522 304866 706758
rect 305102 706522 364546 706758
rect 364782 706522 364866 706758
rect 365102 706522 424546 706758
rect 424782 706522 424866 706758
rect 425102 706522 484546 706758
rect 484782 706522 484866 706758
rect 485102 706522 544546 706758
rect 544782 706522 544866 706758
rect 545102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 4546 706438
rect 4782 706202 4866 706438
rect 5102 706202 64546 706438
rect 64782 706202 64866 706438
rect 65102 706202 124546 706438
rect 124782 706202 124866 706438
rect 125102 706202 184546 706438
rect 184782 706202 184866 706438
rect 185102 706202 244546 706438
rect 244782 706202 244866 706438
rect 245102 706202 304546 706438
rect 304782 706202 304866 706438
rect 305102 706202 364546 706438
rect 364782 706202 364866 706438
rect 365102 706202 424546 706438
rect 424782 706202 424866 706438
rect 425102 706202 484546 706438
rect 484782 706202 484866 706438
rect 485102 706202 544546 706438
rect 544782 706202 544866 706438
rect 545102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 30826 705798
rect 31062 705562 31146 705798
rect 31382 705562 90826 705798
rect 91062 705562 91146 705798
rect 91382 705562 150826 705798
rect 151062 705562 151146 705798
rect 151382 705562 210826 705798
rect 211062 705562 211146 705798
rect 211382 705562 270826 705798
rect 271062 705562 271146 705798
rect 271382 705562 330826 705798
rect 331062 705562 331146 705798
rect 331382 705562 390826 705798
rect 391062 705562 391146 705798
rect 391382 705562 450826 705798
rect 451062 705562 451146 705798
rect 451382 705562 510826 705798
rect 511062 705562 511146 705798
rect 511382 705562 570826 705798
rect 571062 705562 571146 705798
rect 571382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 30826 705478
rect 31062 705242 31146 705478
rect 31382 705242 90826 705478
rect 91062 705242 91146 705478
rect 91382 705242 150826 705478
rect 151062 705242 151146 705478
rect 151382 705242 210826 705478
rect 211062 705242 211146 705478
rect 211382 705242 270826 705478
rect 271062 705242 271146 705478
rect 271382 705242 330826 705478
rect 331062 705242 331146 705478
rect 331382 705242 390826 705478
rect 391062 705242 391146 705478
rect 391382 705242 450826 705478
rect 451062 705242 451146 705478
rect 451382 705242 510826 705478
rect 511062 705242 511146 705478
rect 511382 705242 570826 705478
rect 571062 705242 571146 705478
rect 571382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 826 704838
rect 1062 704602 1146 704838
rect 1382 704602 60826 704838
rect 61062 704602 61146 704838
rect 61382 704602 120826 704838
rect 121062 704602 121146 704838
rect 121382 704602 180826 704838
rect 181062 704602 181146 704838
rect 181382 704602 240826 704838
rect 241062 704602 241146 704838
rect 241382 704602 300826 704838
rect 301062 704602 301146 704838
rect 301382 704602 360826 704838
rect 361062 704602 361146 704838
rect 361382 704602 420826 704838
rect 421062 704602 421146 704838
rect 421382 704602 480826 704838
rect 481062 704602 481146 704838
rect 481382 704602 540826 704838
rect 541062 704602 541146 704838
rect 541382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 826 704518
rect 1062 704282 1146 704518
rect 1382 704282 60826 704518
rect 61062 704282 61146 704518
rect 61382 704282 120826 704518
rect 121062 704282 121146 704518
rect 121382 704282 180826 704518
rect 181062 704282 181146 704518
rect 181382 704282 240826 704518
rect 241062 704282 241146 704518
rect 241382 704282 300826 704518
rect 301062 704282 301146 704518
rect 301382 704282 360826 704518
rect 361062 704282 361146 704518
rect 361382 704282 420826 704518
rect 421062 704282 421146 704518
rect 421382 704282 480826 704518
rect 481062 704282 481146 704518
rect 481382 704282 540826 704518
rect 541062 704282 541146 704518
rect 541382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -6806 699894 590730 699926
rect -6806 699658 -6774 699894
rect -6538 699658 -6454 699894
rect -6218 699658 38266 699894
rect 38502 699658 38586 699894
rect 38822 699658 98266 699894
rect 98502 699658 98586 699894
rect 98822 699658 158266 699894
rect 158502 699658 158586 699894
rect 158822 699658 218266 699894
rect 218502 699658 218586 699894
rect 218822 699658 278266 699894
rect 278502 699658 278586 699894
rect 278822 699658 338266 699894
rect 338502 699658 338586 699894
rect 338822 699658 398266 699894
rect 398502 699658 398586 699894
rect 398822 699658 458266 699894
rect 458502 699658 458586 699894
rect 458822 699658 518266 699894
rect 518502 699658 518586 699894
rect 518822 699658 578266 699894
rect 578502 699658 578586 699894
rect 578822 699658 590142 699894
rect 590378 699658 590462 699894
rect 590698 699658 590730 699894
rect -6806 699574 590730 699658
rect -6806 699338 -6774 699574
rect -6538 699338 -6454 699574
rect -6218 699338 38266 699574
rect 38502 699338 38586 699574
rect 38822 699338 98266 699574
rect 98502 699338 98586 699574
rect 98822 699338 158266 699574
rect 158502 699338 158586 699574
rect 158822 699338 218266 699574
rect 218502 699338 218586 699574
rect 218822 699338 278266 699574
rect 278502 699338 278586 699574
rect 278822 699338 338266 699574
rect 338502 699338 338586 699574
rect 338822 699338 398266 699574
rect 398502 699338 398586 699574
rect 398822 699338 458266 699574
rect 458502 699338 458586 699574
rect 458822 699338 518266 699574
rect 518502 699338 518586 699574
rect 518822 699338 578266 699574
rect 578502 699338 578586 699574
rect 578822 699338 590142 699574
rect 590378 699338 590462 699574
rect 590698 699338 590730 699574
rect -6806 699306 590730 699338
rect -4886 696174 588810 696206
rect -4886 695938 -4854 696174
rect -4618 695938 -4534 696174
rect -4298 695938 34546 696174
rect 34782 695938 34866 696174
rect 35102 695938 94546 696174
rect 94782 695938 94866 696174
rect 95102 695938 154546 696174
rect 154782 695938 154866 696174
rect 155102 695938 214546 696174
rect 214782 695938 214866 696174
rect 215102 695938 274546 696174
rect 274782 695938 274866 696174
rect 275102 695938 334546 696174
rect 334782 695938 334866 696174
rect 335102 695938 394546 696174
rect 394782 695938 394866 696174
rect 395102 695938 454546 696174
rect 454782 695938 454866 696174
rect 455102 695938 514546 696174
rect 514782 695938 514866 696174
rect 515102 695938 574546 696174
rect 574782 695938 574866 696174
rect 575102 695938 588222 696174
rect 588458 695938 588542 696174
rect 588778 695938 588810 696174
rect -4886 695854 588810 695938
rect -4886 695618 -4854 695854
rect -4618 695618 -4534 695854
rect -4298 695618 34546 695854
rect 34782 695618 34866 695854
rect 35102 695618 94546 695854
rect 94782 695618 94866 695854
rect 95102 695618 154546 695854
rect 154782 695618 154866 695854
rect 155102 695618 214546 695854
rect 214782 695618 214866 695854
rect 215102 695618 274546 695854
rect 274782 695618 274866 695854
rect 275102 695618 334546 695854
rect 334782 695618 334866 695854
rect 335102 695618 394546 695854
rect 394782 695618 394866 695854
rect 395102 695618 454546 695854
rect 454782 695618 454866 695854
rect 455102 695618 514546 695854
rect 514782 695618 514866 695854
rect 515102 695618 574546 695854
rect 574782 695618 574866 695854
rect 575102 695618 588222 695854
rect 588458 695618 588542 695854
rect 588778 695618 588810 695854
rect -4886 695586 588810 695618
rect -2966 692454 586890 692486
rect -2966 692218 -2934 692454
rect -2698 692218 -2614 692454
rect -2378 692218 30826 692454
rect 31062 692218 31146 692454
rect 31382 692218 90826 692454
rect 91062 692218 91146 692454
rect 91382 692218 150826 692454
rect 151062 692218 151146 692454
rect 151382 692218 210826 692454
rect 211062 692218 211146 692454
rect 211382 692218 270826 692454
rect 271062 692218 271146 692454
rect 271382 692218 330826 692454
rect 331062 692218 331146 692454
rect 331382 692218 390826 692454
rect 391062 692218 391146 692454
rect 391382 692218 450826 692454
rect 451062 692218 451146 692454
rect 451382 692218 510826 692454
rect 511062 692218 511146 692454
rect 511382 692218 570826 692454
rect 571062 692218 571146 692454
rect 571382 692218 586302 692454
rect 586538 692218 586622 692454
rect 586858 692218 586890 692454
rect -2966 692134 586890 692218
rect -2966 691898 -2934 692134
rect -2698 691898 -2614 692134
rect -2378 691898 30826 692134
rect 31062 691898 31146 692134
rect 31382 691898 90826 692134
rect 91062 691898 91146 692134
rect 91382 691898 150826 692134
rect 151062 691898 151146 692134
rect 151382 691898 210826 692134
rect 211062 691898 211146 692134
rect 211382 691898 270826 692134
rect 271062 691898 271146 692134
rect 271382 691898 330826 692134
rect 331062 691898 331146 692134
rect 331382 691898 390826 692134
rect 391062 691898 391146 692134
rect 391382 691898 450826 692134
rect 451062 691898 451146 692134
rect 451382 691898 510826 692134
rect 511062 691898 511146 692134
rect 511382 691898 570826 692134
rect 571062 691898 571146 692134
rect 571382 691898 586302 692134
rect 586538 691898 586622 692134
rect 586858 691898 586890 692134
rect -2966 691866 586890 691898
rect -8726 673614 592650 673646
rect -8726 673378 -7734 673614
rect -7498 673378 -7414 673614
rect -7178 673378 11986 673614
rect 12222 673378 12306 673614
rect 12542 673378 71986 673614
rect 72222 673378 72306 673614
rect 72542 673378 131986 673614
rect 132222 673378 132306 673614
rect 132542 673378 191986 673614
rect 192222 673378 192306 673614
rect 192542 673378 251986 673614
rect 252222 673378 252306 673614
rect 252542 673378 311986 673614
rect 312222 673378 312306 673614
rect 312542 673378 371986 673614
rect 372222 673378 372306 673614
rect 372542 673378 431986 673614
rect 432222 673378 432306 673614
rect 432542 673378 491986 673614
rect 492222 673378 492306 673614
rect 492542 673378 551986 673614
rect 552222 673378 552306 673614
rect 552542 673378 591102 673614
rect 591338 673378 591422 673614
rect 591658 673378 592650 673614
rect -8726 673294 592650 673378
rect -8726 673058 -7734 673294
rect -7498 673058 -7414 673294
rect -7178 673058 11986 673294
rect 12222 673058 12306 673294
rect 12542 673058 71986 673294
rect 72222 673058 72306 673294
rect 72542 673058 131986 673294
rect 132222 673058 132306 673294
rect 132542 673058 191986 673294
rect 192222 673058 192306 673294
rect 192542 673058 251986 673294
rect 252222 673058 252306 673294
rect 252542 673058 311986 673294
rect 312222 673058 312306 673294
rect 312542 673058 371986 673294
rect 372222 673058 372306 673294
rect 372542 673058 431986 673294
rect 432222 673058 432306 673294
rect 432542 673058 491986 673294
rect 492222 673058 492306 673294
rect 492542 673058 551986 673294
rect 552222 673058 552306 673294
rect 552542 673058 591102 673294
rect 591338 673058 591422 673294
rect 591658 673058 592650 673294
rect -8726 673026 592650 673058
rect -6806 669894 590730 669926
rect -6806 669658 -5814 669894
rect -5578 669658 -5494 669894
rect -5258 669658 8266 669894
rect 8502 669658 8586 669894
rect 8822 669658 68266 669894
rect 68502 669658 68586 669894
rect 68822 669658 128266 669894
rect 128502 669658 128586 669894
rect 128822 669658 188266 669894
rect 188502 669658 188586 669894
rect 188822 669658 248266 669894
rect 248502 669658 248586 669894
rect 248822 669658 308266 669894
rect 308502 669658 308586 669894
rect 308822 669658 368266 669894
rect 368502 669658 368586 669894
rect 368822 669658 428266 669894
rect 428502 669658 428586 669894
rect 428822 669658 488266 669894
rect 488502 669658 488586 669894
rect 488822 669658 548266 669894
rect 548502 669658 548586 669894
rect 548822 669658 589182 669894
rect 589418 669658 589502 669894
rect 589738 669658 590730 669894
rect -6806 669574 590730 669658
rect -6806 669338 -5814 669574
rect -5578 669338 -5494 669574
rect -5258 669338 8266 669574
rect 8502 669338 8586 669574
rect 8822 669338 68266 669574
rect 68502 669338 68586 669574
rect 68822 669338 128266 669574
rect 128502 669338 128586 669574
rect 128822 669338 188266 669574
rect 188502 669338 188586 669574
rect 188822 669338 248266 669574
rect 248502 669338 248586 669574
rect 248822 669338 308266 669574
rect 308502 669338 308586 669574
rect 308822 669338 368266 669574
rect 368502 669338 368586 669574
rect 368822 669338 428266 669574
rect 428502 669338 428586 669574
rect 428822 669338 488266 669574
rect 488502 669338 488586 669574
rect 488822 669338 548266 669574
rect 548502 669338 548586 669574
rect 548822 669338 589182 669574
rect 589418 669338 589502 669574
rect 589738 669338 590730 669574
rect -6806 669306 590730 669338
rect -4886 666174 588810 666206
rect -4886 665938 -3894 666174
rect -3658 665938 -3574 666174
rect -3338 665938 4546 666174
rect 4782 665938 4866 666174
rect 5102 665938 64546 666174
rect 64782 665938 64866 666174
rect 65102 665938 124546 666174
rect 124782 665938 124866 666174
rect 125102 665938 184546 666174
rect 184782 665938 184866 666174
rect 185102 665938 244546 666174
rect 244782 665938 244866 666174
rect 245102 665938 304546 666174
rect 304782 665938 304866 666174
rect 305102 665938 364546 666174
rect 364782 665938 364866 666174
rect 365102 665938 424546 666174
rect 424782 665938 424866 666174
rect 425102 665938 484546 666174
rect 484782 665938 484866 666174
rect 485102 665938 544546 666174
rect 544782 665938 544866 666174
rect 545102 665938 587262 666174
rect 587498 665938 587582 666174
rect 587818 665938 588810 666174
rect -4886 665854 588810 665938
rect -4886 665618 -3894 665854
rect -3658 665618 -3574 665854
rect -3338 665618 4546 665854
rect 4782 665618 4866 665854
rect 5102 665618 64546 665854
rect 64782 665618 64866 665854
rect 65102 665618 124546 665854
rect 124782 665618 124866 665854
rect 125102 665618 184546 665854
rect 184782 665618 184866 665854
rect 185102 665618 244546 665854
rect 244782 665618 244866 665854
rect 245102 665618 304546 665854
rect 304782 665618 304866 665854
rect 305102 665618 364546 665854
rect 364782 665618 364866 665854
rect 365102 665618 424546 665854
rect 424782 665618 424866 665854
rect 425102 665618 484546 665854
rect 484782 665618 484866 665854
rect 485102 665618 544546 665854
rect 544782 665618 544866 665854
rect 545102 665618 587262 665854
rect 587498 665618 587582 665854
rect 587818 665618 588810 665854
rect -4886 665586 588810 665618
rect -2966 662454 586890 662486
rect -2966 662218 -1974 662454
rect -1738 662218 -1654 662454
rect -1418 662218 826 662454
rect 1062 662218 1146 662454
rect 1382 662218 60826 662454
rect 61062 662218 61146 662454
rect 61382 662218 120826 662454
rect 121062 662218 121146 662454
rect 121382 662218 180826 662454
rect 181062 662218 181146 662454
rect 181382 662218 240826 662454
rect 241062 662218 241146 662454
rect 241382 662218 300826 662454
rect 301062 662218 301146 662454
rect 301382 662218 360826 662454
rect 361062 662218 361146 662454
rect 361382 662218 420826 662454
rect 421062 662218 421146 662454
rect 421382 662218 480826 662454
rect 481062 662218 481146 662454
rect 481382 662218 540826 662454
rect 541062 662218 541146 662454
rect 541382 662218 585342 662454
rect 585578 662218 585662 662454
rect 585898 662218 586890 662454
rect -2966 662134 586890 662218
rect -2966 661898 -1974 662134
rect -1738 661898 -1654 662134
rect -1418 661898 826 662134
rect 1062 661898 1146 662134
rect 1382 661898 60826 662134
rect 61062 661898 61146 662134
rect 61382 661898 120826 662134
rect 121062 661898 121146 662134
rect 121382 661898 180826 662134
rect 181062 661898 181146 662134
rect 181382 661898 240826 662134
rect 241062 661898 241146 662134
rect 241382 661898 300826 662134
rect 301062 661898 301146 662134
rect 301382 661898 360826 662134
rect 361062 661898 361146 662134
rect 361382 661898 420826 662134
rect 421062 661898 421146 662134
rect 421382 661898 480826 662134
rect 481062 661898 481146 662134
rect 481382 661898 540826 662134
rect 541062 661898 541146 662134
rect 541382 661898 585342 662134
rect 585578 661898 585662 662134
rect 585898 661898 586890 662134
rect -2966 661866 586890 661898
rect -8726 643614 592650 643646
rect -8726 643378 -8694 643614
rect -8458 643378 -8374 643614
rect -8138 643378 41986 643614
rect 42222 643378 42306 643614
rect 42542 643378 101986 643614
rect 102222 643378 102306 643614
rect 102542 643378 161986 643614
rect 162222 643378 162306 643614
rect 162542 643378 221986 643614
rect 222222 643378 222306 643614
rect 222542 643378 281986 643614
rect 282222 643378 282306 643614
rect 282542 643378 341986 643614
rect 342222 643378 342306 643614
rect 342542 643378 401986 643614
rect 402222 643378 402306 643614
rect 402542 643378 461986 643614
rect 462222 643378 462306 643614
rect 462542 643378 521986 643614
rect 522222 643378 522306 643614
rect 522542 643378 592062 643614
rect 592298 643378 592382 643614
rect 592618 643378 592650 643614
rect -8726 643294 592650 643378
rect -8726 643058 -8694 643294
rect -8458 643058 -8374 643294
rect -8138 643058 41986 643294
rect 42222 643058 42306 643294
rect 42542 643058 101986 643294
rect 102222 643058 102306 643294
rect 102542 643058 161986 643294
rect 162222 643058 162306 643294
rect 162542 643058 221986 643294
rect 222222 643058 222306 643294
rect 222542 643058 281986 643294
rect 282222 643058 282306 643294
rect 282542 643058 341986 643294
rect 342222 643058 342306 643294
rect 342542 643058 401986 643294
rect 402222 643058 402306 643294
rect 402542 643058 461986 643294
rect 462222 643058 462306 643294
rect 462542 643058 521986 643294
rect 522222 643058 522306 643294
rect 522542 643058 592062 643294
rect 592298 643058 592382 643294
rect 592618 643058 592650 643294
rect -8726 643026 592650 643058
rect -6806 639894 590730 639926
rect -6806 639658 -6774 639894
rect -6538 639658 -6454 639894
rect -6218 639658 38266 639894
rect 38502 639658 38586 639894
rect 38822 639658 98266 639894
rect 98502 639658 98586 639894
rect 98822 639658 158266 639894
rect 158502 639658 158586 639894
rect 158822 639658 218266 639894
rect 218502 639658 218586 639894
rect 218822 639658 278266 639894
rect 278502 639658 278586 639894
rect 278822 639658 338266 639894
rect 338502 639658 338586 639894
rect 338822 639658 398266 639894
rect 398502 639658 398586 639894
rect 398822 639658 458266 639894
rect 458502 639658 458586 639894
rect 458822 639658 518266 639894
rect 518502 639658 518586 639894
rect 518822 639658 578266 639894
rect 578502 639658 578586 639894
rect 578822 639658 590142 639894
rect 590378 639658 590462 639894
rect 590698 639658 590730 639894
rect -6806 639574 590730 639658
rect -6806 639338 -6774 639574
rect -6538 639338 -6454 639574
rect -6218 639338 38266 639574
rect 38502 639338 38586 639574
rect 38822 639338 98266 639574
rect 98502 639338 98586 639574
rect 98822 639338 158266 639574
rect 158502 639338 158586 639574
rect 158822 639338 218266 639574
rect 218502 639338 218586 639574
rect 218822 639338 278266 639574
rect 278502 639338 278586 639574
rect 278822 639338 338266 639574
rect 338502 639338 338586 639574
rect 338822 639338 398266 639574
rect 398502 639338 398586 639574
rect 398822 639338 458266 639574
rect 458502 639338 458586 639574
rect 458822 639338 518266 639574
rect 518502 639338 518586 639574
rect 518822 639338 578266 639574
rect 578502 639338 578586 639574
rect 578822 639338 590142 639574
rect 590378 639338 590462 639574
rect 590698 639338 590730 639574
rect -6806 639306 590730 639338
rect -4886 636174 588810 636206
rect -4886 635938 -4854 636174
rect -4618 635938 -4534 636174
rect -4298 635938 34546 636174
rect 34782 635938 34866 636174
rect 35102 635938 94546 636174
rect 94782 635938 94866 636174
rect 95102 635938 154546 636174
rect 154782 635938 154866 636174
rect 155102 635938 214546 636174
rect 214782 635938 214866 636174
rect 215102 635938 274546 636174
rect 274782 635938 274866 636174
rect 275102 635938 334546 636174
rect 334782 635938 334866 636174
rect 335102 635938 394546 636174
rect 394782 635938 394866 636174
rect 395102 635938 454546 636174
rect 454782 635938 454866 636174
rect 455102 635938 514546 636174
rect 514782 635938 514866 636174
rect 515102 635938 574546 636174
rect 574782 635938 574866 636174
rect 575102 635938 588222 636174
rect 588458 635938 588542 636174
rect 588778 635938 588810 636174
rect -4886 635854 588810 635938
rect -4886 635618 -4854 635854
rect -4618 635618 -4534 635854
rect -4298 635618 34546 635854
rect 34782 635618 34866 635854
rect 35102 635618 94546 635854
rect 94782 635618 94866 635854
rect 95102 635618 154546 635854
rect 154782 635618 154866 635854
rect 155102 635618 214546 635854
rect 214782 635618 214866 635854
rect 215102 635618 274546 635854
rect 274782 635618 274866 635854
rect 275102 635618 334546 635854
rect 334782 635618 334866 635854
rect 335102 635618 394546 635854
rect 394782 635618 394866 635854
rect 395102 635618 454546 635854
rect 454782 635618 454866 635854
rect 455102 635618 514546 635854
rect 514782 635618 514866 635854
rect 515102 635618 574546 635854
rect 574782 635618 574866 635854
rect 575102 635618 588222 635854
rect 588458 635618 588542 635854
rect 588778 635618 588810 635854
rect -4886 635586 588810 635618
rect -2966 632454 586890 632486
rect -2966 632218 -2934 632454
rect -2698 632218 -2614 632454
rect -2378 632218 30826 632454
rect 31062 632218 31146 632454
rect 31382 632218 90826 632454
rect 91062 632218 91146 632454
rect 91382 632218 150826 632454
rect 151062 632218 151146 632454
rect 151382 632218 210826 632454
rect 211062 632218 211146 632454
rect 211382 632218 270826 632454
rect 271062 632218 271146 632454
rect 271382 632218 330826 632454
rect 331062 632218 331146 632454
rect 331382 632218 390826 632454
rect 391062 632218 391146 632454
rect 391382 632218 450826 632454
rect 451062 632218 451146 632454
rect 451382 632218 510826 632454
rect 511062 632218 511146 632454
rect 511382 632218 570826 632454
rect 571062 632218 571146 632454
rect 571382 632218 586302 632454
rect 586538 632218 586622 632454
rect 586858 632218 586890 632454
rect -2966 632134 586890 632218
rect -2966 631898 -2934 632134
rect -2698 631898 -2614 632134
rect -2378 631898 30826 632134
rect 31062 631898 31146 632134
rect 31382 631898 90826 632134
rect 91062 631898 91146 632134
rect 91382 631898 150826 632134
rect 151062 631898 151146 632134
rect 151382 631898 210826 632134
rect 211062 631898 211146 632134
rect 211382 631898 270826 632134
rect 271062 631898 271146 632134
rect 271382 631898 330826 632134
rect 331062 631898 331146 632134
rect 331382 631898 390826 632134
rect 391062 631898 391146 632134
rect 391382 631898 450826 632134
rect 451062 631898 451146 632134
rect 451382 631898 510826 632134
rect 511062 631898 511146 632134
rect 511382 631898 570826 632134
rect 571062 631898 571146 632134
rect 571382 631898 586302 632134
rect 586538 631898 586622 632134
rect 586858 631898 586890 632134
rect -2966 631866 586890 631898
rect -8726 613614 592650 613646
rect -8726 613378 -7734 613614
rect -7498 613378 -7414 613614
rect -7178 613378 11986 613614
rect 12222 613378 12306 613614
rect 12542 613378 71986 613614
rect 72222 613378 72306 613614
rect 72542 613378 131986 613614
rect 132222 613378 132306 613614
rect 132542 613378 191986 613614
rect 192222 613378 192306 613614
rect 192542 613378 251986 613614
rect 252222 613378 252306 613614
rect 252542 613378 311986 613614
rect 312222 613378 312306 613614
rect 312542 613378 371986 613614
rect 372222 613378 372306 613614
rect 372542 613378 431986 613614
rect 432222 613378 432306 613614
rect 432542 613378 491986 613614
rect 492222 613378 492306 613614
rect 492542 613378 551986 613614
rect 552222 613378 552306 613614
rect 552542 613378 591102 613614
rect 591338 613378 591422 613614
rect 591658 613378 592650 613614
rect -8726 613294 592650 613378
rect -8726 613058 -7734 613294
rect -7498 613058 -7414 613294
rect -7178 613058 11986 613294
rect 12222 613058 12306 613294
rect 12542 613058 71986 613294
rect 72222 613058 72306 613294
rect 72542 613058 131986 613294
rect 132222 613058 132306 613294
rect 132542 613058 191986 613294
rect 192222 613058 192306 613294
rect 192542 613058 251986 613294
rect 252222 613058 252306 613294
rect 252542 613058 311986 613294
rect 312222 613058 312306 613294
rect 312542 613058 371986 613294
rect 372222 613058 372306 613294
rect 372542 613058 431986 613294
rect 432222 613058 432306 613294
rect 432542 613058 491986 613294
rect 492222 613058 492306 613294
rect 492542 613058 551986 613294
rect 552222 613058 552306 613294
rect 552542 613058 591102 613294
rect 591338 613058 591422 613294
rect 591658 613058 592650 613294
rect -8726 613026 592650 613058
rect -6806 609894 590730 609926
rect -6806 609658 -5814 609894
rect -5578 609658 -5494 609894
rect -5258 609658 8266 609894
rect 8502 609658 8586 609894
rect 8822 609658 68266 609894
rect 68502 609658 68586 609894
rect 68822 609658 128266 609894
rect 128502 609658 128586 609894
rect 128822 609658 188266 609894
rect 188502 609658 188586 609894
rect 188822 609658 248266 609894
rect 248502 609658 248586 609894
rect 248822 609658 308266 609894
rect 308502 609658 308586 609894
rect 308822 609658 368266 609894
rect 368502 609658 368586 609894
rect 368822 609658 428266 609894
rect 428502 609658 428586 609894
rect 428822 609658 488266 609894
rect 488502 609658 488586 609894
rect 488822 609658 548266 609894
rect 548502 609658 548586 609894
rect 548822 609658 589182 609894
rect 589418 609658 589502 609894
rect 589738 609658 590730 609894
rect -6806 609574 590730 609658
rect -6806 609338 -5814 609574
rect -5578 609338 -5494 609574
rect -5258 609338 8266 609574
rect 8502 609338 8586 609574
rect 8822 609338 68266 609574
rect 68502 609338 68586 609574
rect 68822 609338 128266 609574
rect 128502 609338 128586 609574
rect 128822 609338 188266 609574
rect 188502 609338 188586 609574
rect 188822 609338 248266 609574
rect 248502 609338 248586 609574
rect 248822 609338 308266 609574
rect 308502 609338 308586 609574
rect 308822 609338 368266 609574
rect 368502 609338 368586 609574
rect 368822 609338 428266 609574
rect 428502 609338 428586 609574
rect 428822 609338 488266 609574
rect 488502 609338 488586 609574
rect 488822 609338 548266 609574
rect 548502 609338 548586 609574
rect 548822 609338 589182 609574
rect 589418 609338 589502 609574
rect 589738 609338 590730 609574
rect -6806 609306 590730 609338
rect -4886 606174 588810 606206
rect -4886 605938 -3894 606174
rect -3658 605938 -3574 606174
rect -3338 605938 4546 606174
rect 4782 605938 4866 606174
rect 5102 605938 64546 606174
rect 64782 605938 64866 606174
rect 65102 605938 124546 606174
rect 124782 605938 124866 606174
rect 125102 605938 184546 606174
rect 184782 605938 184866 606174
rect 185102 605938 244546 606174
rect 244782 605938 244866 606174
rect 245102 605938 304546 606174
rect 304782 605938 304866 606174
rect 305102 605938 364546 606174
rect 364782 605938 364866 606174
rect 365102 605938 424546 606174
rect 424782 605938 424866 606174
rect 425102 605938 484546 606174
rect 484782 605938 484866 606174
rect 485102 605938 544546 606174
rect 544782 605938 544866 606174
rect 545102 605938 587262 606174
rect 587498 605938 587582 606174
rect 587818 605938 588810 606174
rect -4886 605854 588810 605938
rect -4886 605618 -3894 605854
rect -3658 605618 -3574 605854
rect -3338 605618 4546 605854
rect 4782 605618 4866 605854
rect 5102 605618 64546 605854
rect 64782 605618 64866 605854
rect 65102 605618 124546 605854
rect 124782 605618 124866 605854
rect 125102 605618 184546 605854
rect 184782 605618 184866 605854
rect 185102 605618 244546 605854
rect 244782 605618 244866 605854
rect 245102 605618 304546 605854
rect 304782 605618 304866 605854
rect 305102 605618 364546 605854
rect 364782 605618 364866 605854
rect 365102 605618 424546 605854
rect 424782 605618 424866 605854
rect 425102 605618 484546 605854
rect 484782 605618 484866 605854
rect 485102 605618 544546 605854
rect 544782 605618 544866 605854
rect 545102 605618 587262 605854
rect 587498 605618 587582 605854
rect 587818 605618 588810 605854
rect -4886 605586 588810 605618
rect -2966 602454 586890 602486
rect -2966 602218 -1974 602454
rect -1738 602218 -1654 602454
rect -1418 602218 826 602454
rect 1062 602218 1146 602454
rect 1382 602218 60826 602454
rect 61062 602218 61146 602454
rect 61382 602218 120826 602454
rect 121062 602218 121146 602454
rect 121382 602218 180826 602454
rect 181062 602218 181146 602454
rect 181382 602218 240826 602454
rect 241062 602218 241146 602454
rect 241382 602218 300826 602454
rect 301062 602218 301146 602454
rect 301382 602218 360826 602454
rect 361062 602218 361146 602454
rect 361382 602218 420826 602454
rect 421062 602218 421146 602454
rect 421382 602218 480826 602454
rect 481062 602218 481146 602454
rect 481382 602218 540826 602454
rect 541062 602218 541146 602454
rect 541382 602218 585342 602454
rect 585578 602218 585662 602454
rect 585898 602218 586890 602454
rect -2966 602134 586890 602218
rect -2966 601898 -1974 602134
rect -1738 601898 -1654 602134
rect -1418 601898 826 602134
rect 1062 601898 1146 602134
rect 1382 601898 60826 602134
rect 61062 601898 61146 602134
rect 61382 601898 120826 602134
rect 121062 601898 121146 602134
rect 121382 601898 180826 602134
rect 181062 601898 181146 602134
rect 181382 601898 240826 602134
rect 241062 601898 241146 602134
rect 241382 601898 300826 602134
rect 301062 601898 301146 602134
rect 301382 601898 360826 602134
rect 361062 601898 361146 602134
rect 361382 601898 420826 602134
rect 421062 601898 421146 602134
rect 421382 601898 480826 602134
rect 481062 601898 481146 602134
rect 481382 601898 540826 602134
rect 541062 601898 541146 602134
rect 541382 601898 585342 602134
rect 585578 601898 585662 602134
rect 585898 601898 586890 602134
rect -2966 601866 586890 601898
rect -8726 583614 592650 583646
rect -8726 583378 -8694 583614
rect -8458 583378 -8374 583614
rect -8138 583378 41986 583614
rect 42222 583378 42306 583614
rect 42542 583378 101986 583614
rect 102222 583378 102306 583614
rect 102542 583378 161986 583614
rect 162222 583378 162306 583614
rect 162542 583378 221986 583614
rect 222222 583378 222306 583614
rect 222542 583378 281986 583614
rect 282222 583378 282306 583614
rect 282542 583378 341986 583614
rect 342222 583378 342306 583614
rect 342542 583378 401986 583614
rect 402222 583378 402306 583614
rect 402542 583378 461986 583614
rect 462222 583378 462306 583614
rect 462542 583378 521986 583614
rect 522222 583378 522306 583614
rect 522542 583378 592062 583614
rect 592298 583378 592382 583614
rect 592618 583378 592650 583614
rect -8726 583294 592650 583378
rect -8726 583058 -8694 583294
rect -8458 583058 -8374 583294
rect -8138 583058 41986 583294
rect 42222 583058 42306 583294
rect 42542 583058 101986 583294
rect 102222 583058 102306 583294
rect 102542 583058 161986 583294
rect 162222 583058 162306 583294
rect 162542 583058 221986 583294
rect 222222 583058 222306 583294
rect 222542 583058 281986 583294
rect 282222 583058 282306 583294
rect 282542 583058 341986 583294
rect 342222 583058 342306 583294
rect 342542 583058 401986 583294
rect 402222 583058 402306 583294
rect 402542 583058 461986 583294
rect 462222 583058 462306 583294
rect 462542 583058 521986 583294
rect 522222 583058 522306 583294
rect 522542 583058 592062 583294
rect 592298 583058 592382 583294
rect 592618 583058 592650 583294
rect -8726 583026 592650 583058
rect -6806 579894 590730 579926
rect -6806 579658 -6774 579894
rect -6538 579658 -6454 579894
rect -6218 579658 38266 579894
rect 38502 579658 38586 579894
rect 38822 579658 98266 579894
rect 98502 579658 98586 579894
rect 98822 579658 158266 579894
rect 158502 579658 158586 579894
rect 158822 579658 218266 579894
rect 218502 579658 218586 579894
rect 218822 579658 278266 579894
rect 278502 579658 278586 579894
rect 278822 579658 338266 579894
rect 338502 579658 338586 579894
rect 338822 579658 398266 579894
rect 398502 579658 398586 579894
rect 398822 579658 458266 579894
rect 458502 579658 458586 579894
rect 458822 579658 518266 579894
rect 518502 579658 518586 579894
rect 518822 579658 578266 579894
rect 578502 579658 578586 579894
rect 578822 579658 590142 579894
rect 590378 579658 590462 579894
rect 590698 579658 590730 579894
rect -6806 579574 590730 579658
rect -6806 579338 -6774 579574
rect -6538 579338 -6454 579574
rect -6218 579338 38266 579574
rect 38502 579338 38586 579574
rect 38822 579338 98266 579574
rect 98502 579338 98586 579574
rect 98822 579338 158266 579574
rect 158502 579338 158586 579574
rect 158822 579338 218266 579574
rect 218502 579338 218586 579574
rect 218822 579338 278266 579574
rect 278502 579338 278586 579574
rect 278822 579338 338266 579574
rect 338502 579338 338586 579574
rect 338822 579338 398266 579574
rect 398502 579338 398586 579574
rect 398822 579338 458266 579574
rect 458502 579338 458586 579574
rect 458822 579338 518266 579574
rect 518502 579338 518586 579574
rect 518822 579338 578266 579574
rect 578502 579338 578586 579574
rect 578822 579338 590142 579574
rect 590378 579338 590462 579574
rect 590698 579338 590730 579574
rect -6806 579306 590730 579338
rect -4886 576174 588810 576206
rect -4886 575938 -4854 576174
rect -4618 575938 -4534 576174
rect -4298 575938 34546 576174
rect 34782 575938 34866 576174
rect 35102 575938 94546 576174
rect 94782 575938 94866 576174
rect 95102 575938 154546 576174
rect 154782 575938 154866 576174
rect 155102 575938 214546 576174
rect 214782 575938 214866 576174
rect 215102 575938 274546 576174
rect 274782 575938 274866 576174
rect 275102 575938 334546 576174
rect 334782 575938 334866 576174
rect 335102 575938 394546 576174
rect 394782 575938 394866 576174
rect 395102 575938 454546 576174
rect 454782 575938 454866 576174
rect 455102 575938 514546 576174
rect 514782 575938 514866 576174
rect 515102 575938 574546 576174
rect 574782 575938 574866 576174
rect 575102 575938 588222 576174
rect 588458 575938 588542 576174
rect 588778 575938 588810 576174
rect -4886 575854 588810 575938
rect -4886 575618 -4854 575854
rect -4618 575618 -4534 575854
rect -4298 575618 34546 575854
rect 34782 575618 34866 575854
rect 35102 575618 94546 575854
rect 94782 575618 94866 575854
rect 95102 575618 154546 575854
rect 154782 575618 154866 575854
rect 155102 575618 214546 575854
rect 214782 575618 214866 575854
rect 215102 575618 274546 575854
rect 274782 575618 274866 575854
rect 275102 575618 334546 575854
rect 334782 575618 334866 575854
rect 335102 575618 394546 575854
rect 394782 575618 394866 575854
rect 395102 575618 454546 575854
rect 454782 575618 454866 575854
rect 455102 575618 514546 575854
rect 514782 575618 514866 575854
rect 515102 575618 574546 575854
rect 574782 575618 574866 575854
rect 575102 575618 588222 575854
rect 588458 575618 588542 575854
rect 588778 575618 588810 575854
rect -4886 575586 588810 575618
rect -2966 572454 586890 572486
rect -2966 572218 -2934 572454
rect -2698 572218 -2614 572454
rect -2378 572218 30826 572454
rect 31062 572218 31146 572454
rect 31382 572218 90826 572454
rect 91062 572218 91146 572454
rect 91382 572218 150826 572454
rect 151062 572218 151146 572454
rect 151382 572218 210826 572454
rect 211062 572218 211146 572454
rect 211382 572218 270826 572454
rect 271062 572218 271146 572454
rect 271382 572218 330826 572454
rect 331062 572218 331146 572454
rect 331382 572218 390826 572454
rect 391062 572218 391146 572454
rect 391382 572218 450826 572454
rect 451062 572218 451146 572454
rect 451382 572218 510826 572454
rect 511062 572218 511146 572454
rect 511382 572218 570826 572454
rect 571062 572218 571146 572454
rect 571382 572218 586302 572454
rect 586538 572218 586622 572454
rect 586858 572218 586890 572454
rect -2966 572134 586890 572218
rect -2966 571898 -2934 572134
rect -2698 571898 -2614 572134
rect -2378 571898 30826 572134
rect 31062 571898 31146 572134
rect 31382 571898 90826 572134
rect 91062 571898 91146 572134
rect 91382 571898 150826 572134
rect 151062 571898 151146 572134
rect 151382 571898 210826 572134
rect 211062 571898 211146 572134
rect 211382 571898 270826 572134
rect 271062 571898 271146 572134
rect 271382 571898 330826 572134
rect 331062 571898 331146 572134
rect 331382 571898 390826 572134
rect 391062 571898 391146 572134
rect 391382 571898 450826 572134
rect 451062 571898 451146 572134
rect 451382 571898 510826 572134
rect 511062 571898 511146 572134
rect 511382 571898 570826 572134
rect 571062 571898 571146 572134
rect 571382 571898 586302 572134
rect 586538 571898 586622 572134
rect 586858 571898 586890 572134
rect -2966 571866 586890 571898
rect -8726 553614 592650 553646
rect -8726 553378 -7734 553614
rect -7498 553378 -7414 553614
rect -7178 553378 11986 553614
rect 12222 553378 12306 553614
rect 12542 553378 71986 553614
rect 72222 553378 72306 553614
rect 72542 553378 131986 553614
rect 132222 553378 132306 553614
rect 132542 553378 191986 553614
rect 192222 553378 192306 553614
rect 192542 553378 251986 553614
rect 252222 553378 252306 553614
rect 252542 553378 311986 553614
rect 312222 553378 312306 553614
rect 312542 553378 371986 553614
rect 372222 553378 372306 553614
rect 372542 553378 431986 553614
rect 432222 553378 432306 553614
rect 432542 553378 491986 553614
rect 492222 553378 492306 553614
rect 492542 553378 551986 553614
rect 552222 553378 552306 553614
rect 552542 553378 591102 553614
rect 591338 553378 591422 553614
rect 591658 553378 592650 553614
rect -8726 553294 592650 553378
rect -8726 553058 -7734 553294
rect -7498 553058 -7414 553294
rect -7178 553058 11986 553294
rect 12222 553058 12306 553294
rect 12542 553058 71986 553294
rect 72222 553058 72306 553294
rect 72542 553058 131986 553294
rect 132222 553058 132306 553294
rect 132542 553058 191986 553294
rect 192222 553058 192306 553294
rect 192542 553058 251986 553294
rect 252222 553058 252306 553294
rect 252542 553058 311986 553294
rect 312222 553058 312306 553294
rect 312542 553058 371986 553294
rect 372222 553058 372306 553294
rect 372542 553058 431986 553294
rect 432222 553058 432306 553294
rect 432542 553058 491986 553294
rect 492222 553058 492306 553294
rect 492542 553058 551986 553294
rect 552222 553058 552306 553294
rect 552542 553058 591102 553294
rect 591338 553058 591422 553294
rect 591658 553058 592650 553294
rect -8726 553026 592650 553058
rect -6806 549894 590730 549926
rect -6806 549658 -5814 549894
rect -5578 549658 -5494 549894
rect -5258 549658 8266 549894
rect 8502 549658 8586 549894
rect 8822 549658 68266 549894
rect 68502 549658 68586 549894
rect 68822 549658 128266 549894
rect 128502 549658 128586 549894
rect 128822 549658 188266 549894
rect 188502 549658 188586 549894
rect 188822 549658 248266 549894
rect 248502 549658 248586 549894
rect 248822 549658 308266 549894
rect 308502 549658 308586 549894
rect 308822 549658 368266 549894
rect 368502 549658 368586 549894
rect 368822 549658 428266 549894
rect 428502 549658 428586 549894
rect 428822 549658 488266 549894
rect 488502 549658 488586 549894
rect 488822 549658 548266 549894
rect 548502 549658 548586 549894
rect 548822 549658 589182 549894
rect 589418 549658 589502 549894
rect 589738 549658 590730 549894
rect -6806 549574 590730 549658
rect -6806 549338 -5814 549574
rect -5578 549338 -5494 549574
rect -5258 549338 8266 549574
rect 8502 549338 8586 549574
rect 8822 549338 68266 549574
rect 68502 549338 68586 549574
rect 68822 549338 128266 549574
rect 128502 549338 128586 549574
rect 128822 549338 188266 549574
rect 188502 549338 188586 549574
rect 188822 549338 248266 549574
rect 248502 549338 248586 549574
rect 248822 549338 308266 549574
rect 308502 549338 308586 549574
rect 308822 549338 368266 549574
rect 368502 549338 368586 549574
rect 368822 549338 428266 549574
rect 428502 549338 428586 549574
rect 428822 549338 488266 549574
rect 488502 549338 488586 549574
rect 488822 549338 548266 549574
rect 548502 549338 548586 549574
rect 548822 549338 589182 549574
rect 589418 549338 589502 549574
rect 589738 549338 590730 549574
rect -6806 549306 590730 549338
rect -4886 546174 588810 546206
rect -4886 545938 -3894 546174
rect -3658 545938 -3574 546174
rect -3338 545938 4546 546174
rect 4782 545938 4866 546174
rect 5102 545938 64546 546174
rect 64782 545938 64866 546174
rect 65102 545938 124546 546174
rect 124782 545938 124866 546174
rect 125102 545938 184546 546174
rect 184782 545938 184866 546174
rect 185102 545938 244546 546174
rect 244782 545938 244866 546174
rect 245102 545938 304546 546174
rect 304782 545938 304866 546174
rect 305102 545938 364546 546174
rect 364782 545938 364866 546174
rect 365102 545938 424546 546174
rect 424782 545938 424866 546174
rect 425102 545938 484546 546174
rect 484782 545938 484866 546174
rect 485102 545938 544546 546174
rect 544782 545938 544866 546174
rect 545102 545938 587262 546174
rect 587498 545938 587582 546174
rect 587818 545938 588810 546174
rect -4886 545854 588810 545938
rect -4886 545618 -3894 545854
rect -3658 545618 -3574 545854
rect -3338 545618 4546 545854
rect 4782 545618 4866 545854
rect 5102 545618 64546 545854
rect 64782 545618 64866 545854
rect 65102 545618 124546 545854
rect 124782 545618 124866 545854
rect 125102 545618 184546 545854
rect 184782 545618 184866 545854
rect 185102 545618 244546 545854
rect 244782 545618 244866 545854
rect 245102 545618 304546 545854
rect 304782 545618 304866 545854
rect 305102 545618 364546 545854
rect 364782 545618 364866 545854
rect 365102 545618 424546 545854
rect 424782 545618 424866 545854
rect 425102 545618 484546 545854
rect 484782 545618 484866 545854
rect 485102 545618 544546 545854
rect 544782 545618 544866 545854
rect 545102 545618 587262 545854
rect 587498 545618 587582 545854
rect 587818 545618 588810 545854
rect -4886 545586 588810 545618
rect -2966 542454 586890 542486
rect -2966 542218 -1974 542454
rect -1738 542218 -1654 542454
rect -1418 542218 826 542454
rect 1062 542218 1146 542454
rect 1382 542218 60826 542454
rect 61062 542218 61146 542454
rect 61382 542218 120826 542454
rect 121062 542218 121146 542454
rect 121382 542218 180826 542454
rect 181062 542218 181146 542454
rect 181382 542218 240826 542454
rect 241062 542218 241146 542454
rect 241382 542218 300826 542454
rect 301062 542218 301146 542454
rect 301382 542218 360826 542454
rect 361062 542218 361146 542454
rect 361382 542218 420826 542454
rect 421062 542218 421146 542454
rect 421382 542218 480826 542454
rect 481062 542218 481146 542454
rect 481382 542218 540826 542454
rect 541062 542218 541146 542454
rect 541382 542218 585342 542454
rect 585578 542218 585662 542454
rect 585898 542218 586890 542454
rect -2966 542134 586890 542218
rect -2966 541898 -1974 542134
rect -1738 541898 -1654 542134
rect -1418 541898 826 542134
rect 1062 541898 1146 542134
rect 1382 541898 60826 542134
rect 61062 541898 61146 542134
rect 61382 541898 120826 542134
rect 121062 541898 121146 542134
rect 121382 541898 180826 542134
rect 181062 541898 181146 542134
rect 181382 541898 240826 542134
rect 241062 541898 241146 542134
rect 241382 541898 300826 542134
rect 301062 541898 301146 542134
rect 301382 541898 360826 542134
rect 361062 541898 361146 542134
rect 361382 541898 420826 542134
rect 421062 541898 421146 542134
rect 421382 541898 480826 542134
rect 481062 541898 481146 542134
rect 481382 541898 540826 542134
rect 541062 541898 541146 542134
rect 541382 541898 585342 542134
rect 585578 541898 585662 542134
rect 585898 541898 586890 542134
rect -2966 541866 586890 541898
rect -8726 523614 592650 523646
rect -8726 523378 -8694 523614
rect -8458 523378 -8374 523614
rect -8138 523378 41986 523614
rect 42222 523378 42306 523614
rect 42542 523378 101986 523614
rect 102222 523378 102306 523614
rect 102542 523378 161986 523614
rect 162222 523378 162306 523614
rect 162542 523378 221986 523614
rect 222222 523378 222306 523614
rect 222542 523378 281986 523614
rect 282222 523378 282306 523614
rect 282542 523378 341986 523614
rect 342222 523378 342306 523614
rect 342542 523378 401986 523614
rect 402222 523378 402306 523614
rect 402542 523378 461986 523614
rect 462222 523378 462306 523614
rect 462542 523378 521986 523614
rect 522222 523378 522306 523614
rect 522542 523378 592062 523614
rect 592298 523378 592382 523614
rect 592618 523378 592650 523614
rect -8726 523294 592650 523378
rect -8726 523058 -8694 523294
rect -8458 523058 -8374 523294
rect -8138 523058 41986 523294
rect 42222 523058 42306 523294
rect 42542 523058 101986 523294
rect 102222 523058 102306 523294
rect 102542 523058 161986 523294
rect 162222 523058 162306 523294
rect 162542 523058 221986 523294
rect 222222 523058 222306 523294
rect 222542 523058 281986 523294
rect 282222 523058 282306 523294
rect 282542 523058 341986 523294
rect 342222 523058 342306 523294
rect 342542 523058 401986 523294
rect 402222 523058 402306 523294
rect 402542 523058 461986 523294
rect 462222 523058 462306 523294
rect 462542 523058 521986 523294
rect 522222 523058 522306 523294
rect 522542 523058 592062 523294
rect 592298 523058 592382 523294
rect 592618 523058 592650 523294
rect -8726 523026 592650 523058
rect -6806 519894 590730 519926
rect -6806 519658 -6774 519894
rect -6538 519658 -6454 519894
rect -6218 519658 38266 519894
rect 38502 519658 38586 519894
rect 38822 519658 98266 519894
rect 98502 519658 98586 519894
rect 98822 519658 158266 519894
rect 158502 519658 158586 519894
rect 158822 519658 218266 519894
rect 218502 519658 218586 519894
rect 218822 519658 278266 519894
rect 278502 519658 278586 519894
rect 278822 519658 338266 519894
rect 338502 519658 338586 519894
rect 338822 519658 398266 519894
rect 398502 519658 398586 519894
rect 398822 519658 458266 519894
rect 458502 519658 458586 519894
rect 458822 519658 518266 519894
rect 518502 519658 518586 519894
rect 518822 519658 578266 519894
rect 578502 519658 578586 519894
rect 578822 519658 590142 519894
rect 590378 519658 590462 519894
rect 590698 519658 590730 519894
rect -6806 519574 590730 519658
rect -6806 519338 -6774 519574
rect -6538 519338 -6454 519574
rect -6218 519338 38266 519574
rect 38502 519338 38586 519574
rect 38822 519338 98266 519574
rect 98502 519338 98586 519574
rect 98822 519338 158266 519574
rect 158502 519338 158586 519574
rect 158822 519338 218266 519574
rect 218502 519338 218586 519574
rect 218822 519338 278266 519574
rect 278502 519338 278586 519574
rect 278822 519338 338266 519574
rect 338502 519338 338586 519574
rect 338822 519338 398266 519574
rect 398502 519338 398586 519574
rect 398822 519338 458266 519574
rect 458502 519338 458586 519574
rect 458822 519338 518266 519574
rect 518502 519338 518586 519574
rect 518822 519338 578266 519574
rect 578502 519338 578586 519574
rect 578822 519338 590142 519574
rect 590378 519338 590462 519574
rect 590698 519338 590730 519574
rect -6806 519306 590730 519338
rect -4886 516174 588810 516206
rect -4886 515938 -4854 516174
rect -4618 515938 -4534 516174
rect -4298 515938 34546 516174
rect 34782 515938 34866 516174
rect 35102 515938 94546 516174
rect 94782 515938 94866 516174
rect 95102 515938 154546 516174
rect 154782 515938 154866 516174
rect 155102 515938 214546 516174
rect 214782 515938 214866 516174
rect 215102 515938 274546 516174
rect 274782 515938 274866 516174
rect 275102 515938 334546 516174
rect 334782 515938 334866 516174
rect 335102 515938 394546 516174
rect 394782 515938 394866 516174
rect 395102 515938 454546 516174
rect 454782 515938 454866 516174
rect 455102 515938 514546 516174
rect 514782 515938 514866 516174
rect 515102 515938 574546 516174
rect 574782 515938 574866 516174
rect 575102 515938 588222 516174
rect 588458 515938 588542 516174
rect 588778 515938 588810 516174
rect -4886 515854 588810 515938
rect -4886 515618 -4854 515854
rect -4618 515618 -4534 515854
rect -4298 515618 34546 515854
rect 34782 515618 34866 515854
rect 35102 515618 94546 515854
rect 94782 515618 94866 515854
rect 95102 515618 154546 515854
rect 154782 515618 154866 515854
rect 155102 515618 214546 515854
rect 214782 515618 214866 515854
rect 215102 515618 274546 515854
rect 274782 515618 274866 515854
rect 275102 515618 334546 515854
rect 334782 515618 334866 515854
rect 335102 515618 394546 515854
rect 394782 515618 394866 515854
rect 395102 515618 454546 515854
rect 454782 515618 454866 515854
rect 455102 515618 514546 515854
rect 514782 515618 514866 515854
rect 515102 515618 574546 515854
rect 574782 515618 574866 515854
rect 575102 515618 588222 515854
rect 588458 515618 588542 515854
rect 588778 515618 588810 515854
rect -4886 515586 588810 515618
rect -2966 512454 586890 512486
rect -2966 512218 -2934 512454
rect -2698 512218 -2614 512454
rect -2378 512218 30826 512454
rect 31062 512218 31146 512454
rect 31382 512218 90826 512454
rect 91062 512218 91146 512454
rect 91382 512218 150826 512454
rect 151062 512218 151146 512454
rect 151382 512218 210826 512454
rect 211062 512218 211146 512454
rect 211382 512218 270826 512454
rect 271062 512218 271146 512454
rect 271382 512218 330826 512454
rect 331062 512218 331146 512454
rect 331382 512218 390826 512454
rect 391062 512218 391146 512454
rect 391382 512218 450826 512454
rect 451062 512218 451146 512454
rect 451382 512218 510826 512454
rect 511062 512218 511146 512454
rect 511382 512218 570826 512454
rect 571062 512218 571146 512454
rect 571382 512218 586302 512454
rect 586538 512218 586622 512454
rect 586858 512218 586890 512454
rect -2966 512134 586890 512218
rect -2966 511898 -2934 512134
rect -2698 511898 -2614 512134
rect -2378 511898 30826 512134
rect 31062 511898 31146 512134
rect 31382 511898 90826 512134
rect 91062 511898 91146 512134
rect 91382 511898 150826 512134
rect 151062 511898 151146 512134
rect 151382 511898 210826 512134
rect 211062 511898 211146 512134
rect 211382 511898 270826 512134
rect 271062 511898 271146 512134
rect 271382 511898 330826 512134
rect 331062 511898 331146 512134
rect 331382 511898 390826 512134
rect 391062 511898 391146 512134
rect 391382 511898 450826 512134
rect 451062 511898 451146 512134
rect 451382 511898 510826 512134
rect 511062 511898 511146 512134
rect 511382 511898 570826 512134
rect 571062 511898 571146 512134
rect 571382 511898 586302 512134
rect 586538 511898 586622 512134
rect 586858 511898 586890 512134
rect -2966 511866 586890 511898
rect -8726 493614 592650 493646
rect -8726 493378 -7734 493614
rect -7498 493378 -7414 493614
rect -7178 493378 11986 493614
rect 12222 493378 12306 493614
rect 12542 493378 71986 493614
rect 72222 493378 72306 493614
rect 72542 493378 131986 493614
rect 132222 493378 132306 493614
rect 132542 493378 191986 493614
rect 192222 493378 192306 493614
rect 192542 493378 251986 493614
rect 252222 493378 252306 493614
rect 252542 493378 311986 493614
rect 312222 493378 312306 493614
rect 312542 493378 371986 493614
rect 372222 493378 372306 493614
rect 372542 493378 431986 493614
rect 432222 493378 432306 493614
rect 432542 493378 491986 493614
rect 492222 493378 492306 493614
rect 492542 493378 551986 493614
rect 552222 493378 552306 493614
rect 552542 493378 591102 493614
rect 591338 493378 591422 493614
rect 591658 493378 592650 493614
rect -8726 493294 592650 493378
rect -8726 493058 -7734 493294
rect -7498 493058 -7414 493294
rect -7178 493058 11986 493294
rect 12222 493058 12306 493294
rect 12542 493058 71986 493294
rect 72222 493058 72306 493294
rect 72542 493058 131986 493294
rect 132222 493058 132306 493294
rect 132542 493058 191986 493294
rect 192222 493058 192306 493294
rect 192542 493058 251986 493294
rect 252222 493058 252306 493294
rect 252542 493058 311986 493294
rect 312222 493058 312306 493294
rect 312542 493058 371986 493294
rect 372222 493058 372306 493294
rect 372542 493058 431986 493294
rect 432222 493058 432306 493294
rect 432542 493058 491986 493294
rect 492222 493058 492306 493294
rect 492542 493058 551986 493294
rect 552222 493058 552306 493294
rect 552542 493058 591102 493294
rect 591338 493058 591422 493294
rect 591658 493058 592650 493294
rect -8726 493026 592650 493058
rect -6806 489894 590730 489926
rect -6806 489658 -5814 489894
rect -5578 489658 -5494 489894
rect -5258 489658 8266 489894
rect 8502 489658 8586 489894
rect 8822 489658 68266 489894
rect 68502 489658 68586 489894
rect 68822 489658 128266 489894
rect 128502 489658 128586 489894
rect 128822 489658 188266 489894
rect 188502 489658 188586 489894
rect 188822 489658 248266 489894
rect 248502 489658 248586 489894
rect 248822 489658 308266 489894
rect 308502 489658 308586 489894
rect 308822 489658 368266 489894
rect 368502 489658 368586 489894
rect 368822 489658 428266 489894
rect 428502 489658 428586 489894
rect 428822 489658 488266 489894
rect 488502 489658 488586 489894
rect 488822 489658 548266 489894
rect 548502 489658 548586 489894
rect 548822 489658 589182 489894
rect 589418 489658 589502 489894
rect 589738 489658 590730 489894
rect -6806 489574 590730 489658
rect -6806 489338 -5814 489574
rect -5578 489338 -5494 489574
rect -5258 489338 8266 489574
rect 8502 489338 8586 489574
rect 8822 489338 68266 489574
rect 68502 489338 68586 489574
rect 68822 489338 128266 489574
rect 128502 489338 128586 489574
rect 128822 489338 188266 489574
rect 188502 489338 188586 489574
rect 188822 489338 248266 489574
rect 248502 489338 248586 489574
rect 248822 489338 308266 489574
rect 308502 489338 308586 489574
rect 308822 489338 368266 489574
rect 368502 489338 368586 489574
rect 368822 489338 428266 489574
rect 428502 489338 428586 489574
rect 428822 489338 488266 489574
rect 488502 489338 488586 489574
rect 488822 489338 548266 489574
rect 548502 489338 548586 489574
rect 548822 489338 589182 489574
rect 589418 489338 589502 489574
rect 589738 489338 590730 489574
rect -6806 489306 590730 489338
rect -4886 486174 588810 486206
rect -4886 485938 -3894 486174
rect -3658 485938 -3574 486174
rect -3338 485938 4546 486174
rect 4782 485938 4866 486174
rect 5102 485938 64546 486174
rect 64782 485938 64866 486174
rect 65102 485938 124546 486174
rect 124782 485938 124866 486174
rect 125102 485938 184546 486174
rect 184782 485938 184866 486174
rect 185102 485938 244546 486174
rect 244782 485938 244866 486174
rect 245102 485938 304546 486174
rect 304782 485938 304866 486174
rect 305102 485938 364546 486174
rect 364782 485938 364866 486174
rect 365102 485938 424546 486174
rect 424782 485938 424866 486174
rect 425102 485938 484546 486174
rect 484782 485938 484866 486174
rect 485102 485938 544546 486174
rect 544782 485938 544866 486174
rect 545102 485938 587262 486174
rect 587498 485938 587582 486174
rect 587818 485938 588810 486174
rect -4886 485854 588810 485938
rect -4886 485618 -3894 485854
rect -3658 485618 -3574 485854
rect -3338 485618 4546 485854
rect 4782 485618 4866 485854
rect 5102 485618 64546 485854
rect 64782 485618 64866 485854
rect 65102 485618 124546 485854
rect 124782 485618 124866 485854
rect 125102 485618 184546 485854
rect 184782 485618 184866 485854
rect 185102 485618 244546 485854
rect 244782 485618 244866 485854
rect 245102 485618 304546 485854
rect 304782 485618 304866 485854
rect 305102 485618 364546 485854
rect 364782 485618 364866 485854
rect 365102 485618 424546 485854
rect 424782 485618 424866 485854
rect 425102 485618 484546 485854
rect 484782 485618 484866 485854
rect 485102 485618 544546 485854
rect 544782 485618 544866 485854
rect 545102 485618 587262 485854
rect 587498 485618 587582 485854
rect 587818 485618 588810 485854
rect -4886 485586 588810 485618
rect -2966 482454 586890 482486
rect -2966 482218 -1974 482454
rect -1738 482218 -1654 482454
rect -1418 482218 826 482454
rect 1062 482218 1146 482454
rect 1382 482218 60826 482454
rect 61062 482218 61146 482454
rect 61382 482218 120826 482454
rect 121062 482218 121146 482454
rect 121382 482218 180826 482454
rect 181062 482218 181146 482454
rect 181382 482218 240826 482454
rect 241062 482218 241146 482454
rect 241382 482218 300826 482454
rect 301062 482218 301146 482454
rect 301382 482218 360826 482454
rect 361062 482218 361146 482454
rect 361382 482218 420826 482454
rect 421062 482218 421146 482454
rect 421382 482218 480826 482454
rect 481062 482218 481146 482454
rect 481382 482218 540826 482454
rect 541062 482218 541146 482454
rect 541382 482218 585342 482454
rect 585578 482218 585662 482454
rect 585898 482218 586890 482454
rect -2966 482134 586890 482218
rect -2966 481898 -1974 482134
rect -1738 481898 -1654 482134
rect -1418 481898 826 482134
rect 1062 481898 1146 482134
rect 1382 481898 60826 482134
rect 61062 481898 61146 482134
rect 61382 481898 120826 482134
rect 121062 481898 121146 482134
rect 121382 481898 180826 482134
rect 181062 481898 181146 482134
rect 181382 481898 240826 482134
rect 241062 481898 241146 482134
rect 241382 481898 300826 482134
rect 301062 481898 301146 482134
rect 301382 481898 360826 482134
rect 361062 481898 361146 482134
rect 361382 481898 420826 482134
rect 421062 481898 421146 482134
rect 421382 481898 480826 482134
rect 481062 481898 481146 482134
rect 481382 481898 540826 482134
rect 541062 481898 541146 482134
rect 541382 481898 585342 482134
rect 585578 481898 585662 482134
rect 585898 481898 586890 482134
rect -2966 481866 586890 481898
rect -8726 463614 592650 463646
rect -8726 463378 -8694 463614
rect -8458 463378 -8374 463614
rect -8138 463378 41986 463614
rect 42222 463378 42306 463614
rect 42542 463378 101986 463614
rect 102222 463378 102306 463614
rect 102542 463378 161986 463614
rect 162222 463378 162306 463614
rect 162542 463378 221986 463614
rect 222222 463378 222306 463614
rect 222542 463378 281986 463614
rect 282222 463378 282306 463614
rect 282542 463378 341986 463614
rect 342222 463378 342306 463614
rect 342542 463378 401986 463614
rect 402222 463378 402306 463614
rect 402542 463378 461986 463614
rect 462222 463378 462306 463614
rect 462542 463378 521986 463614
rect 522222 463378 522306 463614
rect 522542 463378 592062 463614
rect 592298 463378 592382 463614
rect 592618 463378 592650 463614
rect -8726 463294 592650 463378
rect -8726 463058 -8694 463294
rect -8458 463058 -8374 463294
rect -8138 463058 41986 463294
rect 42222 463058 42306 463294
rect 42542 463058 101986 463294
rect 102222 463058 102306 463294
rect 102542 463058 161986 463294
rect 162222 463058 162306 463294
rect 162542 463058 221986 463294
rect 222222 463058 222306 463294
rect 222542 463058 281986 463294
rect 282222 463058 282306 463294
rect 282542 463058 341986 463294
rect 342222 463058 342306 463294
rect 342542 463058 401986 463294
rect 402222 463058 402306 463294
rect 402542 463058 461986 463294
rect 462222 463058 462306 463294
rect 462542 463058 521986 463294
rect 522222 463058 522306 463294
rect 522542 463058 592062 463294
rect 592298 463058 592382 463294
rect 592618 463058 592650 463294
rect -8726 463026 592650 463058
rect -6806 459894 590730 459926
rect -6806 459658 -6774 459894
rect -6538 459658 -6454 459894
rect -6218 459658 38266 459894
rect 38502 459658 38586 459894
rect 38822 459658 98266 459894
rect 98502 459658 98586 459894
rect 98822 459658 158266 459894
rect 158502 459658 158586 459894
rect 158822 459658 218266 459894
rect 218502 459658 218586 459894
rect 218822 459658 278266 459894
rect 278502 459658 278586 459894
rect 278822 459658 338266 459894
rect 338502 459658 338586 459894
rect 338822 459658 398266 459894
rect 398502 459658 398586 459894
rect 398822 459658 458266 459894
rect 458502 459658 458586 459894
rect 458822 459658 518266 459894
rect 518502 459658 518586 459894
rect 518822 459658 578266 459894
rect 578502 459658 578586 459894
rect 578822 459658 590142 459894
rect 590378 459658 590462 459894
rect 590698 459658 590730 459894
rect -6806 459574 590730 459658
rect -6806 459338 -6774 459574
rect -6538 459338 -6454 459574
rect -6218 459338 38266 459574
rect 38502 459338 38586 459574
rect 38822 459338 98266 459574
rect 98502 459338 98586 459574
rect 98822 459338 158266 459574
rect 158502 459338 158586 459574
rect 158822 459338 218266 459574
rect 218502 459338 218586 459574
rect 218822 459338 278266 459574
rect 278502 459338 278586 459574
rect 278822 459338 338266 459574
rect 338502 459338 338586 459574
rect 338822 459338 398266 459574
rect 398502 459338 398586 459574
rect 398822 459338 458266 459574
rect 458502 459338 458586 459574
rect 458822 459338 518266 459574
rect 518502 459338 518586 459574
rect 518822 459338 578266 459574
rect 578502 459338 578586 459574
rect 578822 459338 590142 459574
rect 590378 459338 590462 459574
rect 590698 459338 590730 459574
rect -6806 459306 590730 459338
rect -4886 456174 588810 456206
rect -4886 455938 -4854 456174
rect -4618 455938 -4534 456174
rect -4298 455938 34546 456174
rect 34782 455938 34866 456174
rect 35102 455938 94546 456174
rect 94782 455938 94866 456174
rect 95102 455938 154546 456174
rect 154782 455938 154866 456174
rect 155102 455938 214546 456174
rect 214782 455938 214866 456174
rect 215102 455938 274546 456174
rect 274782 455938 274866 456174
rect 275102 455938 334546 456174
rect 334782 455938 334866 456174
rect 335102 455938 394546 456174
rect 394782 455938 394866 456174
rect 395102 455938 454546 456174
rect 454782 455938 454866 456174
rect 455102 455938 514546 456174
rect 514782 455938 514866 456174
rect 515102 455938 574546 456174
rect 574782 455938 574866 456174
rect 575102 455938 588222 456174
rect 588458 455938 588542 456174
rect 588778 455938 588810 456174
rect -4886 455854 588810 455938
rect -4886 455618 -4854 455854
rect -4618 455618 -4534 455854
rect -4298 455618 34546 455854
rect 34782 455618 34866 455854
rect 35102 455618 94546 455854
rect 94782 455618 94866 455854
rect 95102 455618 154546 455854
rect 154782 455618 154866 455854
rect 155102 455618 214546 455854
rect 214782 455618 214866 455854
rect 215102 455618 274546 455854
rect 274782 455618 274866 455854
rect 275102 455618 334546 455854
rect 334782 455618 334866 455854
rect 335102 455618 394546 455854
rect 394782 455618 394866 455854
rect 395102 455618 454546 455854
rect 454782 455618 454866 455854
rect 455102 455618 514546 455854
rect 514782 455618 514866 455854
rect 515102 455618 574546 455854
rect 574782 455618 574866 455854
rect 575102 455618 588222 455854
rect 588458 455618 588542 455854
rect 588778 455618 588810 455854
rect -4886 455586 588810 455618
rect -2966 452454 586890 452486
rect -2966 452218 -2934 452454
rect -2698 452218 -2614 452454
rect -2378 452218 30826 452454
rect 31062 452218 31146 452454
rect 31382 452218 90826 452454
rect 91062 452218 91146 452454
rect 91382 452218 150826 452454
rect 151062 452218 151146 452454
rect 151382 452218 210826 452454
rect 211062 452218 211146 452454
rect 211382 452218 270826 452454
rect 271062 452218 271146 452454
rect 271382 452218 330826 452454
rect 331062 452218 331146 452454
rect 331382 452218 390826 452454
rect 391062 452218 391146 452454
rect 391382 452218 450826 452454
rect 451062 452218 451146 452454
rect 451382 452218 510826 452454
rect 511062 452218 511146 452454
rect 511382 452218 570826 452454
rect 571062 452218 571146 452454
rect 571382 452218 586302 452454
rect 586538 452218 586622 452454
rect 586858 452218 586890 452454
rect -2966 452134 586890 452218
rect -2966 451898 -2934 452134
rect -2698 451898 -2614 452134
rect -2378 451898 30826 452134
rect 31062 451898 31146 452134
rect 31382 451898 90826 452134
rect 91062 451898 91146 452134
rect 91382 451898 150826 452134
rect 151062 451898 151146 452134
rect 151382 451898 210826 452134
rect 211062 451898 211146 452134
rect 211382 451898 270826 452134
rect 271062 451898 271146 452134
rect 271382 451898 330826 452134
rect 331062 451898 331146 452134
rect 331382 451898 390826 452134
rect 391062 451898 391146 452134
rect 391382 451898 450826 452134
rect 451062 451898 451146 452134
rect 451382 451898 510826 452134
rect 511062 451898 511146 452134
rect 511382 451898 570826 452134
rect 571062 451898 571146 452134
rect 571382 451898 586302 452134
rect 586538 451898 586622 452134
rect 586858 451898 586890 452134
rect -2966 451866 586890 451898
rect -8726 433614 592650 433646
rect -8726 433378 -7734 433614
rect -7498 433378 -7414 433614
rect -7178 433378 11986 433614
rect 12222 433378 12306 433614
rect 12542 433378 71986 433614
rect 72222 433378 72306 433614
rect 72542 433378 131986 433614
rect 132222 433378 132306 433614
rect 132542 433378 191986 433614
rect 192222 433378 192306 433614
rect 192542 433378 251986 433614
rect 252222 433378 252306 433614
rect 252542 433378 311986 433614
rect 312222 433378 312306 433614
rect 312542 433378 371986 433614
rect 372222 433378 372306 433614
rect 372542 433378 431986 433614
rect 432222 433378 432306 433614
rect 432542 433378 491986 433614
rect 492222 433378 492306 433614
rect 492542 433378 551986 433614
rect 552222 433378 552306 433614
rect 552542 433378 591102 433614
rect 591338 433378 591422 433614
rect 591658 433378 592650 433614
rect -8726 433294 592650 433378
rect -8726 433058 -7734 433294
rect -7498 433058 -7414 433294
rect -7178 433058 11986 433294
rect 12222 433058 12306 433294
rect 12542 433058 71986 433294
rect 72222 433058 72306 433294
rect 72542 433058 131986 433294
rect 132222 433058 132306 433294
rect 132542 433058 191986 433294
rect 192222 433058 192306 433294
rect 192542 433058 251986 433294
rect 252222 433058 252306 433294
rect 252542 433058 311986 433294
rect 312222 433058 312306 433294
rect 312542 433058 371986 433294
rect 372222 433058 372306 433294
rect 372542 433058 431986 433294
rect 432222 433058 432306 433294
rect 432542 433058 491986 433294
rect 492222 433058 492306 433294
rect 492542 433058 551986 433294
rect 552222 433058 552306 433294
rect 552542 433058 591102 433294
rect 591338 433058 591422 433294
rect 591658 433058 592650 433294
rect -8726 433026 592650 433058
rect -6806 429894 590730 429926
rect -6806 429658 -5814 429894
rect -5578 429658 -5494 429894
rect -5258 429658 8266 429894
rect 8502 429658 8586 429894
rect 8822 429658 68266 429894
rect 68502 429658 68586 429894
rect 68822 429658 128266 429894
rect 128502 429658 128586 429894
rect 128822 429658 188266 429894
rect 188502 429658 188586 429894
rect 188822 429658 248266 429894
rect 248502 429658 248586 429894
rect 248822 429658 308266 429894
rect 308502 429658 308586 429894
rect 308822 429658 368266 429894
rect 368502 429658 368586 429894
rect 368822 429658 428266 429894
rect 428502 429658 428586 429894
rect 428822 429658 488266 429894
rect 488502 429658 488586 429894
rect 488822 429658 548266 429894
rect 548502 429658 548586 429894
rect 548822 429658 589182 429894
rect 589418 429658 589502 429894
rect 589738 429658 590730 429894
rect -6806 429574 590730 429658
rect -6806 429338 -5814 429574
rect -5578 429338 -5494 429574
rect -5258 429338 8266 429574
rect 8502 429338 8586 429574
rect 8822 429338 68266 429574
rect 68502 429338 68586 429574
rect 68822 429338 128266 429574
rect 128502 429338 128586 429574
rect 128822 429338 188266 429574
rect 188502 429338 188586 429574
rect 188822 429338 248266 429574
rect 248502 429338 248586 429574
rect 248822 429338 308266 429574
rect 308502 429338 308586 429574
rect 308822 429338 368266 429574
rect 368502 429338 368586 429574
rect 368822 429338 428266 429574
rect 428502 429338 428586 429574
rect 428822 429338 488266 429574
rect 488502 429338 488586 429574
rect 488822 429338 548266 429574
rect 548502 429338 548586 429574
rect 548822 429338 589182 429574
rect 589418 429338 589502 429574
rect 589738 429338 590730 429574
rect -6806 429306 590730 429338
rect -4886 426174 588810 426206
rect -4886 425938 -3894 426174
rect -3658 425938 -3574 426174
rect -3338 425938 4546 426174
rect 4782 425938 4866 426174
rect 5102 425938 64546 426174
rect 64782 425938 64866 426174
rect 65102 425938 124546 426174
rect 124782 425938 124866 426174
rect 125102 425938 184546 426174
rect 184782 425938 184866 426174
rect 185102 425938 244546 426174
rect 244782 425938 244866 426174
rect 245102 425938 304546 426174
rect 304782 425938 304866 426174
rect 305102 425938 364546 426174
rect 364782 425938 364866 426174
rect 365102 425938 424546 426174
rect 424782 425938 424866 426174
rect 425102 425938 484546 426174
rect 484782 425938 484866 426174
rect 485102 425938 544546 426174
rect 544782 425938 544866 426174
rect 545102 425938 587262 426174
rect 587498 425938 587582 426174
rect 587818 425938 588810 426174
rect -4886 425854 588810 425938
rect -4886 425618 -3894 425854
rect -3658 425618 -3574 425854
rect -3338 425618 4546 425854
rect 4782 425618 4866 425854
rect 5102 425618 64546 425854
rect 64782 425618 64866 425854
rect 65102 425618 124546 425854
rect 124782 425618 124866 425854
rect 125102 425618 184546 425854
rect 184782 425618 184866 425854
rect 185102 425618 244546 425854
rect 244782 425618 244866 425854
rect 245102 425618 304546 425854
rect 304782 425618 304866 425854
rect 305102 425618 364546 425854
rect 364782 425618 364866 425854
rect 365102 425618 424546 425854
rect 424782 425618 424866 425854
rect 425102 425618 484546 425854
rect 484782 425618 484866 425854
rect 485102 425618 544546 425854
rect 544782 425618 544866 425854
rect 545102 425618 587262 425854
rect 587498 425618 587582 425854
rect 587818 425618 588810 425854
rect -4886 425586 588810 425618
rect -2966 422454 586890 422486
rect -2966 422218 -1974 422454
rect -1738 422218 -1654 422454
rect -1418 422218 826 422454
rect 1062 422218 1146 422454
rect 1382 422218 60826 422454
rect 61062 422218 61146 422454
rect 61382 422218 120826 422454
rect 121062 422218 121146 422454
rect 121382 422218 180826 422454
rect 181062 422218 181146 422454
rect 181382 422218 240826 422454
rect 241062 422218 241146 422454
rect 241382 422218 300826 422454
rect 301062 422218 301146 422454
rect 301382 422218 360826 422454
rect 361062 422218 361146 422454
rect 361382 422218 420826 422454
rect 421062 422218 421146 422454
rect 421382 422218 480826 422454
rect 481062 422218 481146 422454
rect 481382 422218 540826 422454
rect 541062 422218 541146 422454
rect 541382 422218 585342 422454
rect 585578 422218 585662 422454
rect 585898 422218 586890 422454
rect -2966 422134 586890 422218
rect -2966 421898 -1974 422134
rect -1738 421898 -1654 422134
rect -1418 421898 826 422134
rect 1062 421898 1146 422134
rect 1382 421898 60826 422134
rect 61062 421898 61146 422134
rect 61382 421898 120826 422134
rect 121062 421898 121146 422134
rect 121382 421898 180826 422134
rect 181062 421898 181146 422134
rect 181382 421898 240826 422134
rect 241062 421898 241146 422134
rect 241382 421898 300826 422134
rect 301062 421898 301146 422134
rect 301382 421898 360826 422134
rect 361062 421898 361146 422134
rect 361382 421898 420826 422134
rect 421062 421898 421146 422134
rect 421382 421898 480826 422134
rect 481062 421898 481146 422134
rect 481382 421898 540826 422134
rect 541062 421898 541146 422134
rect 541382 421898 585342 422134
rect 585578 421898 585662 422134
rect 585898 421898 586890 422134
rect -2966 421866 586890 421898
rect -8726 403614 592650 403646
rect -8726 403378 -8694 403614
rect -8458 403378 -8374 403614
rect -8138 403378 41986 403614
rect 42222 403378 42306 403614
rect 42542 403378 101986 403614
rect 102222 403378 102306 403614
rect 102542 403378 161986 403614
rect 162222 403378 162306 403614
rect 162542 403378 221986 403614
rect 222222 403378 222306 403614
rect 222542 403378 281986 403614
rect 282222 403378 282306 403614
rect 282542 403378 341986 403614
rect 342222 403378 342306 403614
rect 342542 403378 401986 403614
rect 402222 403378 402306 403614
rect 402542 403378 461986 403614
rect 462222 403378 462306 403614
rect 462542 403378 521986 403614
rect 522222 403378 522306 403614
rect 522542 403378 592062 403614
rect 592298 403378 592382 403614
rect 592618 403378 592650 403614
rect -8726 403294 592650 403378
rect -8726 403058 -8694 403294
rect -8458 403058 -8374 403294
rect -8138 403058 41986 403294
rect 42222 403058 42306 403294
rect 42542 403058 101986 403294
rect 102222 403058 102306 403294
rect 102542 403058 161986 403294
rect 162222 403058 162306 403294
rect 162542 403058 221986 403294
rect 222222 403058 222306 403294
rect 222542 403058 281986 403294
rect 282222 403058 282306 403294
rect 282542 403058 341986 403294
rect 342222 403058 342306 403294
rect 342542 403058 401986 403294
rect 402222 403058 402306 403294
rect 402542 403058 461986 403294
rect 462222 403058 462306 403294
rect 462542 403058 521986 403294
rect 522222 403058 522306 403294
rect 522542 403058 592062 403294
rect 592298 403058 592382 403294
rect 592618 403058 592650 403294
rect -8726 403026 592650 403058
rect -6806 399894 590730 399926
rect -6806 399658 -6774 399894
rect -6538 399658 -6454 399894
rect -6218 399658 38266 399894
rect 38502 399658 38586 399894
rect 38822 399658 98266 399894
rect 98502 399658 98586 399894
rect 98822 399658 158266 399894
rect 158502 399658 158586 399894
rect 158822 399658 218266 399894
rect 218502 399658 218586 399894
rect 218822 399658 278266 399894
rect 278502 399658 278586 399894
rect 278822 399658 338266 399894
rect 338502 399658 338586 399894
rect 338822 399658 398266 399894
rect 398502 399658 398586 399894
rect 398822 399658 458266 399894
rect 458502 399658 458586 399894
rect 458822 399658 518266 399894
rect 518502 399658 518586 399894
rect 518822 399658 578266 399894
rect 578502 399658 578586 399894
rect 578822 399658 590142 399894
rect 590378 399658 590462 399894
rect 590698 399658 590730 399894
rect -6806 399574 590730 399658
rect -6806 399338 -6774 399574
rect -6538 399338 -6454 399574
rect -6218 399338 38266 399574
rect 38502 399338 38586 399574
rect 38822 399338 98266 399574
rect 98502 399338 98586 399574
rect 98822 399338 158266 399574
rect 158502 399338 158586 399574
rect 158822 399338 218266 399574
rect 218502 399338 218586 399574
rect 218822 399338 278266 399574
rect 278502 399338 278586 399574
rect 278822 399338 338266 399574
rect 338502 399338 338586 399574
rect 338822 399338 398266 399574
rect 398502 399338 398586 399574
rect 398822 399338 458266 399574
rect 458502 399338 458586 399574
rect 458822 399338 518266 399574
rect 518502 399338 518586 399574
rect 518822 399338 578266 399574
rect 578502 399338 578586 399574
rect 578822 399338 590142 399574
rect 590378 399338 590462 399574
rect 590698 399338 590730 399574
rect -6806 399306 590730 399338
rect -4886 396174 588810 396206
rect -4886 395938 -4854 396174
rect -4618 395938 -4534 396174
rect -4298 395938 34546 396174
rect 34782 395938 34866 396174
rect 35102 395938 94546 396174
rect 94782 395938 94866 396174
rect 95102 395938 154546 396174
rect 154782 395938 154866 396174
rect 155102 395938 214546 396174
rect 214782 395938 214866 396174
rect 215102 395938 274546 396174
rect 274782 395938 274866 396174
rect 275102 395938 334546 396174
rect 334782 395938 334866 396174
rect 335102 395938 394546 396174
rect 394782 395938 394866 396174
rect 395102 395938 454546 396174
rect 454782 395938 454866 396174
rect 455102 395938 514546 396174
rect 514782 395938 514866 396174
rect 515102 395938 574546 396174
rect 574782 395938 574866 396174
rect 575102 395938 588222 396174
rect 588458 395938 588542 396174
rect 588778 395938 588810 396174
rect -4886 395854 588810 395938
rect -4886 395618 -4854 395854
rect -4618 395618 -4534 395854
rect -4298 395618 34546 395854
rect 34782 395618 34866 395854
rect 35102 395618 94546 395854
rect 94782 395618 94866 395854
rect 95102 395618 154546 395854
rect 154782 395618 154866 395854
rect 155102 395618 214546 395854
rect 214782 395618 214866 395854
rect 215102 395618 274546 395854
rect 274782 395618 274866 395854
rect 275102 395618 334546 395854
rect 334782 395618 334866 395854
rect 335102 395618 394546 395854
rect 394782 395618 394866 395854
rect 395102 395618 454546 395854
rect 454782 395618 454866 395854
rect 455102 395618 514546 395854
rect 514782 395618 514866 395854
rect 515102 395618 574546 395854
rect 574782 395618 574866 395854
rect 575102 395618 588222 395854
rect 588458 395618 588542 395854
rect 588778 395618 588810 395854
rect -4886 395586 588810 395618
rect -2966 392454 586890 392486
rect -2966 392218 -2934 392454
rect -2698 392218 -2614 392454
rect -2378 392218 30826 392454
rect 31062 392218 31146 392454
rect 31382 392218 90826 392454
rect 91062 392218 91146 392454
rect 91382 392218 150826 392454
rect 151062 392218 151146 392454
rect 151382 392218 210826 392454
rect 211062 392218 211146 392454
rect 211382 392218 270826 392454
rect 271062 392218 271146 392454
rect 271382 392218 330826 392454
rect 331062 392218 331146 392454
rect 331382 392218 390826 392454
rect 391062 392218 391146 392454
rect 391382 392218 450826 392454
rect 451062 392218 451146 392454
rect 451382 392218 510826 392454
rect 511062 392218 511146 392454
rect 511382 392218 570826 392454
rect 571062 392218 571146 392454
rect 571382 392218 586302 392454
rect 586538 392218 586622 392454
rect 586858 392218 586890 392454
rect -2966 392134 586890 392218
rect -2966 391898 -2934 392134
rect -2698 391898 -2614 392134
rect -2378 391898 30826 392134
rect 31062 391898 31146 392134
rect 31382 391898 90826 392134
rect 91062 391898 91146 392134
rect 91382 391898 150826 392134
rect 151062 391898 151146 392134
rect 151382 391898 210826 392134
rect 211062 391898 211146 392134
rect 211382 391898 270826 392134
rect 271062 391898 271146 392134
rect 271382 391898 330826 392134
rect 331062 391898 331146 392134
rect 331382 391898 390826 392134
rect 391062 391898 391146 392134
rect 391382 391898 450826 392134
rect 451062 391898 451146 392134
rect 451382 391898 510826 392134
rect 511062 391898 511146 392134
rect 511382 391898 570826 392134
rect 571062 391898 571146 392134
rect 571382 391898 586302 392134
rect 586538 391898 586622 392134
rect 586858 391898 586890 392134
rect -2966 391866 586890 391898
rect -8726 373614 592650 373646
rect -8726 373378 -7734 373614
rect -7498 373378 -7414 373614
rect -7178 373378 11986 373614
rect 12222 373378 12306 373614
rect 12542 373378 71986 373614
rect 72222 373378 72306 373614
rect 72542 373378 131986 373614
rect 132222 373378 132306 373614
rect 132542 373378 191986 373614
rect 192222 373378 192306 373614
rect 192542 373378 251986 373614
rect 252222 373378 252306 373614
rect 252542 373378 311986 373614
rect 312222 373378 312306 373614
rect 312542 373378 371986 373614
rect 372222 373378 372306 373614
rect 372542 373378 431986 373614
rect 432222 373378 432306 373614
rect 432542 373378 491986 373614
rect 492222 373378 492306 373614
rect 492542 373378 551986 373614
rect 552222 373378 552306 373614
rect 552542 373378 591102 373614
rect 591338 373378 591422 373614
rect 591658 373378 592650 373614
rect -8726 373294 592650 373378
rect -8726 373058 -7734 373294
rect -7498 373058 -7414 373294
rect -7178 373058 11986 373294
rect 12222 373058 12306 373294
rect 12542 373058 71986 373294
rect 72222 373058 72306 373294
rect 72542 373058 131986 373294
rect 132222 373058 132306 373294
rect 132542 373058 191986 373294
rect 192222 373058 192306 373294
rect 192542 373058 251986 373294
rect 252222 373058 252306 373294
rect 252542 373058 311986 373294
rect 312222 373058 312306 373294
rect 312542 373058 371986 373294
rect 372222 373058 372306 373294
rect 372542 373058 431986 373294
rect 432222 373058 432306 373294
rect 432542 373058 491986 373294
rect 492222 373058 492306 373294
rect 492542 373058 551986 373294
rect 552222 373058 552306 373294
rect 552542 373058 591102 373294
rect 591338 373058 591422 373294
rect 591658 373058 592650 373294
rect -8726 373026 592650 373058
rect -6806 369894 590730 369926
rect -6806 369658 -5814 369894
rect -5578 369658 -5494 369894
rect -5258 369658 8266 369894
rect 8502 369658 8586 369894
rect 8822 369658 68266 369894
rect 68502 369658 68586 369894
rect 68822 369658 128266 369894
rect 128502 369658 128586 369894
rect 128822 369658 188266 369894
rect 188502 369658 188586 369894
rect 188822 369658 248266 369894
rect 248502 369658 248586 369894
rect 248822 369658 308266 369894
rect 308502 369658 308586 369894
rect 308822 369658 368266 369894
rect 368502 369658 368586 369894
rect 368822 369658 428266 369894
rect 428502 369658 428586 369894
rect 428822 369658 488266 369894
rect 488502 369658 488586 369894
rect 488822 369658 548266 369894
rect 548502 369658 548586 369894
rect 548822 369658 589182 369894
rect 589418 369658 589502 369894
rect 589738 369658 590730 369894
rect -6806 369574 590730 369658
rect -6806 369338 -5814 369574
rect -5578 369338 -5494 369574
rect -5258 369338 8266 369574
rect 8502 369338 8586 369574
rect 8822 369338 68266 369574
rect 68502 369338 68586 369574
rect 68822 369338 128266 369574
rect 128502 369338 128586 369574
rect 128822 369338 188266 369574
rect 188502 369338 188586 369574
rect 188822 369338 248266 369574
rect 248502 369338 248586 369574
rect 248822 369338 308266 369574
rect 308502 369338 308586 369574
rect 308822 369338 368266 369574
rect 368502 369338 368586 369574
rect 368822 369338 428266 369574
rect 428502 369338 428586 369574
rect 428822 369338 488266 369574
rect 488502 369338 488586 369574
rect 488822 369338 548266 369574
rect 548502 369338 548586 369574
rect 548822 369338 589182 369574
rect 589418 369338 589502 369574
rect 589738 369338 590730 369574
rect -6806 369306 590730 369338
rect -4886 366174 588810 366206
rect -4886 365938 -3894 366174
rect -3658 365938 -3574 366174
rect -3338 365938 4546 366174
rect 4782 365938 4866 366174
rect 5102 365938 64546 366174
rect 64782 365938 64866 366174
rect 65102 365938 124546 366174
rect 124782 365938 124866 366174
rect 125102 365938 184546 366174
rect 184782 365938 184866 366174
rect 185102 365938 244546 366174
rect 244782 365938 244866 366174
rect 245102 365938 304546 366174
rect 304782 365938 304866 366174
rect 305102 365938 364546 366174
rect 364782 365938 364866 366174
rect 365102 365938 424546 366174
rect 424782 365938 424866 366174
rect 425102 365938 484546 366174
rect 484782 365938 484866 366174
rect 485102 365938 544546 366174
rect 544782 365938 544866 366174
rect 545102 365938 587262 366174
rect 587498 365938 587582 366174
rect 587818 365938 588810 366174
rect -4886 365854 588810 365938
rect -4886 365618 -3894 365854
rect -3658 365618 -3574 365854
rect -3338 365618 4546 365854
rect 4782 365618 4866 365854
rect 5102 365618 64546 365854
rect 64782 365618 64866 365854
rect 65102 365618 124546 365854
rect 124782 365618 124866 365854
rect 125102 365618 184546 365854
rect 184782 365618 184866 365854
rect 185102 365618 244546 365854
rect 244782 365618 244866 365854
rect 245102 365618 304546 365854
rect 304782 365618 304866 365854
rect 305102 365618 364546 365854
rect 364782 365618 364866 365854
rect 365102 365618 424546 365854
rect 424782 365618 424866 365854
rect 425102 365618 484546 365854
rect 484782 365618 484866 365854
rect 485102 365618 544546 365854
rect 544782 365618 544866 365854
rect 545102 365618 587262 365854
rect 587498 365618 587582 365854
rect 587818 365618 588810 365854
rect -4886 365586 588810 365618
rect -2966 362454 586890 362486
rect -2966 362218 -1974 362454
rect -1738 362218 -1654 362454
rect -1418 362218 826 362454
rect 1062 362218 1146 362454
rect 1382 362218 60826 362454
rect 61062 362218 61146 362454
rect 61382 362218 120826 362454
rect 121062 362218 121146 362454
rect 121382 362218 180826 362454
rect 181062 362218 181146 362454
rect 181382 362218 240826 362454
rect 241062 362218 241146 362454
rect 241382 362218 300826 362454
rect 301062 362218 301146 362454
rect 301382 362218 360826 362454
rect 361062 362218 361146 362454
rect 361382 362218 420826 362454
rect 421062 362218 421146 362454
rect 421382 362218 480826 362454
rect 481062 362218 481146 362454
rect 481382 362218 540826 362454
rect 541062 362218 541146 362454
rect 541382 362218 585342 362454
rect 585578 362218 585662 362454
rect 585898 362218 586890 362454
rect -2966 362134 586890 362218
rect -2966 361898 -1974 362134
rect -1738 361898 -1654 362134
rect -1418 361898 826 362134
rect 1062 361898 1146 362134
rect 1382 361898 60826 362134
rect 61062 361898 61146 362134
rect 61382 361898 120826 362134
rect 121062 361898 121146 362134
rect 121382 361898 180826 362134
rect 181062 361898 181146 362134
rect 181382 361898 240826 362134
rect 241062 361898 241146 362134
rect 241382 361898 300826 362134
rect 301062 361898 301146 362134
rect 301382 361898 360826 362134
rect 361062 361898 361146 362134
rect 361382 361898 420826 362134
rect 421062 361898 421146 362134
rect 421382 361898 480826 362134
rect 481062 361898 481146 362134
rect 481382 361898 540826 362134
rect 541062 361898 541146 362134
rect 541382 361898 585342 362134
rect 585578 361898 585662 362134
rect 585898 361898 586890 362134
rect -2966 361866 586890 361898
rect -8726 343614 592650 343646
rect -8726 343378 -8694 343614
rect -8458 343378 -8374 343614
rect -8138 343378 41986 343614
rect 42222 343378 42306 343614
rect 42542 343378 101986 343614
rect 102222 343378 102306 343614
rect 102542 343378 161986 343614
rect 162222 343378 162306 343614
rect 162542 343378 221986 343614
rect 222222 343378 222306 343614
rect 222542 343378 281986 343614
rect 282222 343378 282306 343614
rect 282542 343378 341986 343614
rect 342222 343378 342306 343614
rect 342542 343378 401986 343614
rect 402222 343378 402306 343614
rect 402542 343378 461986 343614
rect 462222 343378 462306 343614
rect 462542 343378 521986 343614
rect 522222 343378 522306 343614
rect 522542 343378 592062 343614
rect 592298 343378 592382 343614
rect 592618 343378 592650 343614
rect -8726 343294 592650 343378
rect -8726 343058 -8694 343294
rect -8458 343058 -8374 343294
rect -8138 343058 41986 343294
rect 42222 343058 42306 343294
rect 42542 343058 101986 343294
rect 102222 343058 102306 343294
rect 102542 343058 161986 343294
rect 162222 343058 162306 343294
rect 162542 343058 221986 343294
rect 222222 343058 222306 343294
rect 222542 343058 281986 343294
rect 282222 343058 282306 343294
rect 282542 343058 341986 343294
rect 342222 343058 342306 343294
rect 342542 343058 401986 343294
rect 402222 343058 402306 343294
rect 402542 343058 461986 343294
rect 462222 343058 462306 343294
rect 462542 343058 521986 343294
rect 522222 343058 522306 343294
rect 522542 343058 592062 343294
rect 592298 343058 592382 343294
rect 592618 343058 592650 343294
rect -8726 343026 592650 343058
rect -6806 339894 590730 339926
rect -6806 339658 -6774 339894
rect -6538 339658 -6454 339894
rect -6218 339658 38266 339894
rect 38502 339658 38586 339894
rect 38822 339658 98266 339894
rect 98502 339658 98586 339894
rect 98822 339658 158266 339894
rect 158502 339658 158586 339894
rect 158822 339658 218266 339894
rect 218502 339658 218586 339894
rect 218822 339658 278266 339894
rect 278502 339658 278586 339894
rect 278822 339658 338266 339894
rect 338502 339658 338586 339894
rect 338822 339658 398266 339894
rect 398502 339658 398586 339894
rect 398822 339658 458266 339894
rect 458502 339658 458586 339894
rect 458822 339658 518266 339894
rect 518502 339658 518586 339894
rect 518822 339658 578266 339894
rect 578502 339658 578586 339894
rect 578822 339658 590142 339894
rect 590378 339658 590462 339894
rect 590698 339658 590730 339894
rect -6806 339574 590730 339658
rect -6806 339338 -6774 339574
rect -6538 339338 -6454 339574
rect -6218 339338 38266 339574
rect 38502 339338 38586 339574
rect 38822 339338 98266 339574
rect 98502 339338 98586 339574
rect 98822 339338 158266 339574
rect 158502 339338 158586 339574
rect 158822 339338 218266 339574
rect 218502 339338 218586 339574
rect 218822 339338 278266 339574
rect 278502 339338 278586 339574
rect 278822 339338 338266 339574
rect 338502 339338 338586 339574
rect 338822 339338 398266 339574
rect 398502 339338 398586 339574
rect 398822 339338 458266 339574
rect 458502 339338 458586 339574
rect 458822 339338 518266 339574
rect 518502 339338 518586 339574
rect 518822 339338 578266 339574
rect 578502 339338 578586 339574
rect 578822 339338 590142 339574
rect 590378 339338 590462 339574
rect 590698 339338 590730 339574
rect -6806 339306 590730 339338
rect -4886 336174 588810 336206
rect -4886 335938 -4854 336174
rect -4618 335938 -4534 336174
rect -4298 335938 34546 336174
rect 34782 335938 34866 336174
rect 35102 335938 94546 336174
rect 94782 335938 94866 336174
rect 95102 335938 154546 336174
rect 154782 335938 154866 336174
rect 155102 335938 214546 336174
rect 214782 335938 214866 336174
rect 215102 335938 274546 336174
rect 274782 335938 274866 336174
rect 275102 335938 334546 336174
rect 334782 335938 334866 336174
rect 335102 335938 394546 336174
rect 394782 335938 394866 336174
rect 395102 335938 454546 336174
rect 454782 335938 454866 336174
rect 455102 335938 514546 336174
rect 514782 335938 514866 336174
rect 515102 335938 574546 336174
rect 574782 335938 574866 336174
rect 575102 335938 588222 336174
rect 588458 335938 588542 336174
rect 588778 335938 588810 336174
rect -4886 335854 588810 335938
rect -4886 335618 -4854 335854
rect -4618 335618 -4534 335854
rect -4298 335618 34546 335854
rect 34782 335618 34866 335854
rect 35102 335618 94546 335854
rect 94782 335618 94866 335854
rect 95102 335618 154546 335854
rect 154782 335618 154866 335854
rect 155102 335618 214546 335854
rect 214782 335618 214866 335854
rect 215102 335618 274546 335854
rect 274782 335618 274866 335854
rect 275102 335618 334546 335854
rect 334782 335618 334866 335854
rect 335102 335618 394546 335854
rect 394782 335618 394866 335854
rect 395102 335618 454546 335854
rect 454782 335618 454866 335854
rect 455102 335618 514546 335854
rect 514782 335618 514866 335854
rect 515102 335618 574546 335854
rect 574782 335618 574866 335854
rect 575102 335618 588222 335854
rect 588458 335618 588542 335854
rect 588778 335618 588810 335854
rect -4886 335586 588810 335618
rect -2966 332454 586890 332486
rect -2966 332218 -2934 332454
rect -2698 332218 -2614 332454
rect -2378 332218 30826 332454
rect 31062 332218 31146 332454
rect 31382 332218 90826 332454
rect 91062 332218 91146 332454
rect 91382 332218 150826 332454
rect 151062 332218 151146 332454
rect 151382 332218 210826 332454
rect 211062 332218 211146 332454
rect 211382 332218 270826 332454
rect 271062 332218 271146 332454
rect 271382 332218 330826 332454
rect 331062 332218 331146 332454
rect 331382 332218 390826 332454
rect 391062 332218 391146 332454
rect 391382 332218 450826 332454
rect 451062 332218 451146 332454
rect 451382 332218 510826 332454
rect 511062 332218 511146 332454
rect 511382 332218 570826 332454
rect 571062 332218 571146 332454
rect 571382 332218 586302 332454
rect 586538 332218 586622 332454
rect 586858 332218 586890 332454
rect -2966 332134 586890 332218
rect -2966 331898 -2934 332134
rect -2698 331898 -2614 332134
rect -2378 331898 30826 332134
rect 31062 331898 31146 332134
rect 31382 331898 90826 332134
rect 91062 331898 91146 332134
rect 91382 331898 150826 332134
rect 151062 331898 151146 332134
rect 151382 331898 210826 332134
rect 211062 331898 211146 332134
rect 211382 331898 270826 332134
rect 271062 331898 271146 332134
rect 271382 331898 330826 332134
rect 331062 331898 331146 332134
rect 331382 331898 390826 332134
rect 391062 331898 391146 332134
rect 391382 331898 450826 332134
rect 451062 331898 451146 332134
rect 451382 331898 510826 332134
rect 511062 331898 511146 332134
rect 511382 331898 570826 332134
rect 571062 331898 571146 332134
rect 571382 331898 586302 332134
rect 586538 331898 586622 332134
rect 586858 331898 586890 332134
rect -2966 331866 586890 331898
rect -8726 313614 592650 313646
rect -8726 313378 -7734 313614
rect -7498 313378 -7414 313614
rect -7178 313378 11986 313614
rect 12222 313378 12306 313614
rect 12542 313378 71986 313614
rect 72222 313378 72306 313614
rect 72542 313378 131986 313614
rect 132222 313378 132306 313614
rect 132542 313378 191986 313614
rect 192222 313378 192306 313614
rect 192542 313378 251986 313614
rect 252222 313378 252306 313614
rect 252542 313378 311986 313614
rect 312222 313378 312306 313614
rect 312542 313378 371986 313614
rect 372222 313378 372306 313614
rect 372542 313378 431986 313614
rect 432222 313378 432306 313614
rect 432542 313378 491986 313614
rect 492222 313378 492306 313614
rect 492542 313378 551986 313614
rect 552222 313378 552306 313614
rect 552542 313378 591102 313614
rect 591338 313378 591422 313614
rect 591658 313378 592650 313614
rect -8726 313294 592650 313378
rect -8726 313058 -7734 313294
rect -7498 313058 -7414 313294
rect -7178 313058 11986 313294
rect 12222 313058 12306 313294
rect 12542 313058 71986 313294
rect 72222 313058 72306 313294
rect 72542 313058 131986 313294
rect 132222 313058 132306 313294
rect 132542 313058 191986 313294
rect 192222 313058 192306 313294
rect 192542 313058 251986 313294
rect 252222 313058 252306 313294
rect 252542 313058 311986 313294
rect 312222 313058 312306 313294
rect 312542 313058 371986 313294
rect 372222 313058 372306 313294
rect 372542 313058 431986 313294
rect 432222 313058 432306 313294
rect 432542 313058 491986 313294
rect 492222 313058 492306 313294
rect 492542 313058 551986 313294
rect 552222 313058 552306 313294
rect 552542 313058 591102 313294
rect 591338 313058 591422 313294
rect 591658 313058 592650 313294
rect -8726 313026 592650 313058
rect -6806 309894 590730 309926
rect -6806 309658 -5814 309894
rect -5578 309658 -5494 309894
rect -5258 309658 8266 309894
rect 8502 309658 8586 309894
rect 8822 309658 68266 309894
rect 68502 309658 68586 309894
rect 68822 309658 128266 309894
rect 128502 309658 128586 309894
rect 128822 309658 188266 309894
rect 188502 309658 188586 309894
rect 188822 309658 248266 309894
rect 248502 309658 248586 309894
rect 248822 309658 308266 309894
rect 308502 309658 308586 309894
rect 308822 309658 368266 309894
rect 368502 309658 368586 309894
rect 368822 309658 428266 309894
rect 428502 309658 428586 309894
rect 428822 309658 488266 309894
rect 488502 309658 488586 309894
rect 488822 309658 548266 309894
rect 548502 309658 548586 309894
rect 548822 309658 589182 309894
rect 589418 309658 589502 309894
rect 589738 309658 590730 309894
rect -6806 309574 590730 309658
rect -6806 309338 -5814 309574
rect -5578 309338 -5494 309574
rect -5258 309338 8266 309574
rect 8502 309338 8586 309574
rect 8822 309338 68266 309574
rect 68502 309338 68586 309574
rect 68822 309338 128266 309574
rect 128502 309338 128586 309574
rect 128822 309338 188266 309574
rect 188502 309338 188586 309574
rect 188822 309338 248266 309574
rect 248502 309338 248586 309574
rect 248822 309338 308266 309574
rect 308502 309338 308586 309574
rect 308822 309338 368266 309574
rect 368502 309338 368586 309574
rect 368822 309338 428266 309574
rect 428502 309338 428586 309574
rect 428822 309338 488266 309574
rect 488502 309338 488586 309574
rect 488822 309338 548266 309574
rect 548502 309338 548586 309574
rect 548822 309338 589182 309574
rect 589418 309338 589502 309574
rect 589738 309338 590730 309574
rect -6806 309306 590730 309338
rect -4886 306174 588810 306206
rect -4886 305938 -3894 306174
rect -3658 305938 -3574 306174
rect -3338 305938 4546 306174
rect 4782 305938 4866 306174
rect 5102 305938 64546 306174
rect 64782 305938 64866 306174
rect 65102 305938 124546 306174
rect 124782 305938 124866 306174
rect 125102 305938 184546 306174
rect 184782 305938 184866 306174
rect 185102 305938 244546 306174
rect 244782 305938 244866 306174
rect 245102 305938 304546 306174
rect 304782 305938 304866 306174
rect 305102 305938 364546 306174
rect 364782 305938 364866 306174
rect 365102 305938 424546 306174
rect 424782 305938 424866 306174
rect 425102 305938 484546 306174
rect 484782 305938 484866 306174
rect 485102 305938 544546 306174
rect 544782 305938 544866 306174
rect 545102 305938 587262 306174
rect 587498 305938 587582 306174
rect 587818 305938 588810 306174
rect -4886 305854 588810 305938
rect -4886 305618 -3894 305854
rect -3658 305618 -3574 305854
rect -3338 305618 4546 305854
rect 4782 305618 4866 305854
rect 5102 305618 64546 305854
rect 64782 305618 64866 305854
rect 65102 305618 124546 305854
rect 124782 305618 124866 305854
rect 125102 305618 184546 305854
rect 184782 305618 184866 305854
rect 185102 305618 244546 305854
rect 244782 305618 244866 305854
rect 245102 305618 304546 305854
rect 304782 305618 304866 305854
rect 305102 305618 364546 305854
rect 364782 305618 364866 305854
rect 365102 305618 424546 305854
rect 424782 305618 424866 305854
rect 425102 305618 484546 305854
rect 484782 305618 484866 305854
rect 485102 305618 544546 305854
rect 544782 305618 544866 305854
rect 545102 305618 587262 305854
rect 587498 305618 587582 305854
rect 587818 305618 588810 305854
rect -4886 305586 588810 305618
rect -2966 302454 586890 302486
rect -2966 302218 -1974 302454
rect -1738 302218 -1654 302454
rect -1418 302218 826 302454
rect 1062 302218 1146 302454
rect 1382 302218 60826 302454
rect 61062 302218 61146 302454
rect 61382 302218 120826 302454
rect 121062 302218 121146 302454
rect 121382 302218 180826 302454
rect 181062 302218 181146 302454
rect 181382 302218 240826 302454
rect 241062 302218 241146 302454
rect 241382 302218 300826 302454
rect 301062 302218 301146 302454
rect 301382 302218 360826 302454
rect 361062 302218 361146 302454
rect 361382 302218 420826 302454
rect 421062 302218 421146 302454
rect 421382 302218 480826 302454
rect 481062 302218 481146 302454
rect 481382 302218 540826 302454
rect 541062 302218 541146 302454
rect 541382 302218 585342 302454
rect 585578 302218 585662 302454
rect 585898 302218 586890 302454
rect -2966 302134 586890 302218
rect -2966 301898 -1974 302134
rect -1738 301898 -1654 302134
rect -1418 301898 826 302134
rect 1062 301898 1146 302134
rect 1382 301898 60826 302134
rect 61062 301898 61146 302134
rect 61382 301898 120826 302134
rect 121062 301898 121146 302134
rect 121382 301898 180826 302134
rect 181062 301898 181146 302134
rect 181382 301898 240826 302134
rect 241062 301898 241146 302134
rect 241382 301898 300826 302134
rect 301062 301898 301146 302134
rect 301382 301898 360826 302134
rect 361062 301898 361146 302134
rect 361382 301898 420826 302134
rect 421062 301898 421146 302134
rect 421382 301898 480826 302134
rect 481062 301898 481146 302134
rect 481382 301898 540826 302134
rect 541062 301898 541146 302134
rect 541382 301898 585342 302134
rect 585578 301898 585662 302134
rect 585898 301898 586890 302134
rect -2966 301866 586890 301898
rect -8726 283614 592650 283646
rect -8726 283378 -8694 283614
rect -8458 283378 -8374 283614
rect -8138 283378 41986 283614
rect 42222 283378 42306 283614
rect 42542 283378 101986 283614
rect 102222 283378 102306 283614
rect 102542 283378 161986 283614
rect 162222 283378 162306 283614
rect 162542 283378 221986 283614
rect 222222 283378 222306 283614
rect 222542 283378 281986 283614
rect 282222 283378 282306 283614
rect 282542 283378 341986 283614
rect 342222 283378 342306 283614
rect 342542 283378 401986 283614
rect 402222 283378 402306 283614
rect 402542 283378 461986 283614
rect 462222 283378 462306 283614
rect 462542 283378 521986 283614
rect 522222 283378 522306 283614
rect 522542 283378 592062 283614
rect 592298 283378 592382 283614
rect 592618 283378 592650 283614
rect -8726 283294 592650 283378
rect -8726 283058 -8694 283294
rect -8458 283058 -8374 283294
rect -8138 283058 41986 283294
rect 42222 283058 42306 283294
rect 42542 283058 101986 283294
rect 102222 283058 102306 283294
rect 102542 283058 161986 283294
rect 162222 283058 162306 283294
rect 162542 283058 221986 283294
rect 222222 283058 222306 283294
rect 222542 283058 281986 283294
rect 282222 283058 282306 283294
rect 282542 283058 341986 283294
rect 342222 283058 342306 283294
rect 342542 283058 401986 283294
rect 402222 283058 402306 283294
rect 402542 283058 461986 283294
rect 462222 283058 462306 283294
rect 462542 283058 521986 283294
rect 522222 283058 522306 283294
rect 522542 283058 592062 283294
rect 592298 283058 592382 283294
rect 592618 283058 592650 283294
rect -8726 283026 592650 283058
rect -6806 279894 590730 279926
rect -6806 279658 -6774 279894
rect -6538 279658 -6454 279894
rect -6218 279658 38266 279894
rect 38502 279658 38586 279894
rect 38822 279658 98266 279894
rect 98502 279658 98586 279894
rect 98822 279658 158266 279894
rect 158502 279658 158586 279894
rect 158822 279658 218266 279894
rect 218502 279658 218586 279894
rect 218822 279658 278266 279894
rect 278502 279658 278586 279894
rect 278822 279658 338266 279894
rect 338502 279658 338586 279894
rect 338822 279658 398266 279894
rect 398502 279658 398586 279894
rect 398822 279658 458266 279894
rect 458502 279658 458586 279894
rect 458822 279658 518266 279894
rect 518502 279658 518586 279894
rect 518822 279658 578266 279894
rect 578502 279658 578586 279894
rect 578822 279658 590142 279894
rect 590378 279658 590462 279894
rect 590698 279658 590730 279894
rect -6806 279574 590730 279658
rect -6806 279338 -6774 279574
rect -6538 279338 -6454 279574
rect -6218 279338 38266 279574
rect 38502 279338 38586 279574
rect 38822 279338 98266 279574
rect 98502 279338 98586 279574
rect 98822 279338 158266 279574
rect 158502 279338 158586 279574
rect 158822 279338 218266 279574
rect 218502 279338 218586 279574
rect 218822 279338 278266 279574
rect 278502 279338 278586 279574
rect 278822 279338 338266 279574
rect 338502 279338 338586 279574
rect 338822 279338 398266 279574
rect 398502 279338 398586 279574
rect 398822 279338 458266 279574
rect 458502 279338 458586 279574
rect 458822 279338 518266 279574
rect 518502 279338 518586 279574
rect 518822 279338 578266 279574
rect 578502 279338 578586 279574
rect 578822 279338 590142 279574
rect 590378 279338 590462 279574
rect 590698 279338 590730 279574
rect -6806 279306 590730 279338
rect -4886 276174 588810 276206
rect -4886 275938 -4854 276174
rect -4618 275938 -4534 276174
rect -4298 275938 34546 276174
rect 34782 275938 34866 276174
rect 35102 275938 94546 276174
rect 94782 275938 94866 276174
rect 95102 275938 154546 276174
rect 154782 275938 154866 276174
rect 155102 275938 214546 276174
rect 214782 275938 214866 276174
rect 215102 275938 274546 276174
rect 274782 275938 274866 276174
rect 275102 275938 334546 276174
rect 334782 275938 334866 276174
rect 335102 275938 394546 276174
rect 394782 275938 394866 276174
rect 395102 275938 454546 276174
rect 454782 275938 454866 276174
rect 455102 275938 514546 276174
rect 514782 275938 514866 276174
rect 515102 275938 574546 276174
rect 574782 275938 574866 276174
rect 575102 275938 588222 276174
rect 588458 275938 588542 276174
rect 588778 275938 588810 276174
rect -4886 275854 588810 275938
rect -4886 275618 -4854 275854
rect -4618 275618 -4534 275854
rect -4298 275618 34546 275854
rect 34782 275618 34866 275854
rect 35102 275618 94546 275854
rect 94782 275618 94866 275854
rect 95102 275618 154546 275854
rect 154782 275618 154866 275854
rect 155102 275618 214546 275854
rect 214782 275618 214866 275854
rect 215102 275618 274546 275854
rect 274782 275618 274866 275854
rect 275102 275618 334546 275854
rect 334782 275618 334866 275854
rect 335102 275618 394546 275854
rect 394782 275618 394866 275854
rect 395102 275618 454546 275854
rect 454782 275618 454866 275854
rect 455102 275618 514546 275854
rect 514782 275618 514866 275854
rect 515102 275618 574546 275854
rect 574782 275618 574866 275854
rect 575102 275618 588222 275854
rect 588458 275618 588542 275854
rect 588778 275618 588810 275854
rect -4886 275586 588810 275618
rect -2966 272454 586890 272486
rect -2966 272218 -2934 272454
rect -2698 272218 -2614 272454
rect -2378 272218 30826 272454
rect 31062 272218 31146 272454
rect 31382 272218 90826 272454
rect 91062 272218 91146 272454
rect 91382 272218 150826 272454
rect 151062 272218 151146 272454
rect 151382 272218 210826 272454
rect 211062 272218 211146 272454
rect 211382 272218 270826 272454
rect 271062 272218 271146 272454
rect 271382 272218 330826 272454
rect 331062 272218 331146 272454
rect 331382 272218 390826 272454
rect 391062 272218 391146 272454
rect 391382 272218 450826 272454
rect 451062 272218 451146 272454
rect 451382 272218 510826 272454
rect 511062 272218 511146 272454
rect 511382 272218 570826 272454
rect 571062 272218 571146 272454
rect 571382 272218 586302 272454
rect 586538 272218 586622 272454
rect 586858 272218 586890 272454
rect -2966 272134 586890 272218
rect -2966 271898 -2934 272134
rect -2698 271898 -2614 272134
rect -2378 271898 30826 272134
rect 31062 271898 31146 272134
rect 31382 271898 90826 272134
rect 91062 271898 91146 272134
rect 91382 271898 150826 272134
rect 151062 271898 151146 272134
rect 151382 271898 210826 272134
rect 211062 271898 211146 272134
rect 211382 271898 270826 272134
rect 271062 271898 271146 272134
rect 271382 271898 330826 272134
rect 331062 271898 331146 272134
rect 331382 271898 390826 272134
rect 391062 271898 391146 272134
rect 391382 271898 450826 272134
rect 451062 271898 451146 272134
rect 451382 271898 510826 272134
rect 511062 271898 511146 272134
rect 511382 271898 570826 272134
rect 571062 271898 571146 272134
rect 571382 271898 586302 272134
rect 586538 271898 586622 272134
rect 586858 271898 586890 272134
rect -2966 271866 586890 271898
rect -8726 253614 592650 253646
rect -8726 253378 -7734 253614
rect -7498 253378 -7414 253614
rect -7178 253378 11986 253614
rect 12222 253378 12306 253614
rect 12542 253378 71986 253614
rect 72222 253378 72306 253614
rect 72542 253378 131986 253614
rect 132222 253378 132306 253614
rect 132542 253378 191986 253614
rect 192222 253378 192306 253614
rect 192542 253378 311986 253614
rect 312222 253378 312306 253614
rect 312542 253378 371986 253614
rect 372222 253378 372306 253614
rect 372542 253378 431986 253614
rect 432222 253378 432306 253614
rect 432542 253378 491986 253614
rect 492222 253378 492306 253614
rect 492542 253378 551986 253614
rect 552222 253378 552306 253614
rect 552542 253378 591102 253614
rect 591338 253378 591422 253614
rect 591658 253378 592650 253614
rect -8726 253294 592650 253378
rect -8726 253058 -7734 253294
rect -7498 253058 -7414 253294
rect -7178 253058 11986 253294
rect 12222 253058 12306 253294
rect 12542 253058 71986 253294
rect 72222 253058 72306 253294
rect 72542 253058 131986 253294
rect 132222 253058 132306 253294
rect 132542 253058 191986 253294
rect 192222 253058 192306 253294
rect 192542 253058 311986 253294
rect 312222 253058 312306 253294
rect 312542 253058 371986 253294
rect 372222 253058 372306 253294
rect 372542 253058 431986 253294
rect 432222 253058 432306 253294
rect 432542 253058 491986 253294
rect 492222 253058 492306 253294
rect 492542 253058 551986 253294
rect 552222 253058 552306 253294
rect 552542 253058 591102 253294
rect 591338 253058 591422 253294
rect 591658 253058 592650 253294
rect -8726 253026 592650 253058
rect -6806 249894 590730 249926
rect -6806 249658 -5814 249894
rect -5578 249658 -5494 249894
rect -5258 249658 8266 249894
rect 8502 249658 8586 249894
rect 8822 249658 68266 249894
rect 68502 249658 68586 249894
rect 68822 249658 128266 249894
rect 128502 249658 128586 249894
rect 128822 249658 188266 249894
rect 188502 249658 188586 249894
rect 188822 249658 308266 249894
rect 308502 249658 308586 249894
rect 308822 249658 368266 249894
rect 368502 249658 368586 249894
rect 368822 249658 428266 249894
rect 428502 249658 428586 249894
rect 428822 249658 488266 249894
rect 488502 249658 488586 249894
rect 488822 249658 548266 249894
rect 548502 249658 548586 249894
rect 548822 249658 589182 249894
rect 589418 249658 589502 249894
rect 589738 249658 590730 249894
rect -6806 249574 590730 249658
rect -6806 249338 -5814 249574
rect -5578 249338 -5494 249574
rect -5258 249338 8266 249574
rect 8502 249338 8586 249574
rect 8822 249338 68266 249574
rect 68502 249338 68586 249574
rect 68822 249338 128266 249574
rect 128502 249338 128586 249574
rect 128822 249338 188266 249574
rect 188502 249338 188586 249574
rect 188822 249338 308266 249574
rect 308502 249338 308586 249574
rect 308822 249338 368266 249574
rect 368502 249338 368586 249574
rect 368822 249338 428266 249574
rect 428502 249338 428586 249574
rect 428822 249338 488266 249574
rect 488502 249338 488586 249574
rect 488822 249338 548266 249574
rect 548502 249338 548586 249574
rect 548822 249338 589182 249574
rect 589418 249338 589502 249574
rect 589738 249338 590730 249574
rect -6806 249306 590730 249338
rect 24588 247298 249756 247340
rect 24588 247062 24630 247298
rect 24866 247062 249478 247298
rect 249714 247062 249756 247298
rect 24588 247020 249756 247062
rect -4886 246174 588810 246206
rect -4886 245938 -3894 246174
rect -3658 245938 -3574 246174
rect -3338 245938 4546 246174
rect 4782 245938 4866 246174
rect 5102 245938 64546 246174
rect 64782 245938 64866 246174
rect 65102 245938 124546 246174
rect 124782 245938 124866 246174
rect 125102 245938 184546 246174
rect 184782 245938 184866 246174
rect 185102 245938 304546 246174
rect 304782 245938 304866 246174
rect 305102 245938 364546 246174
rect 364782 245938 364866 246174
rect 365102 245938 424546 246174
rect 424782 245938 424866 246174
rect 425102 245938 484546 246174
rect 484782 245938 484866 246174
rect 485102 245938 544546 246174
rect 544782 245938 544866 246174
rect 545102 245938 587262 246174
rect 587498 245938 587582 246174
rect 587818 245938 588810 246174
rect -4886 245854 588810 245938
rect -4886 245618 -3894 245854
rect -3658 245618 -3574 245854
rect -3338 245618 4546 245854
rect 4782 245618 4866 245854
rect 5102 245618 64546 245854
rect 64782 245618 64866 245854
rect 65102 245618 124546 245854
rect 124782 245618 124866 245854
rect 125102 245618 184546 245854
rect 184782 245618 184866 245854
rect 185102 245618 304546 245854
rect 304782 245618 304866 245854
rect 305102 245618 364546 245854
rect 364782 245618 364866 245854
rect 365102 245618 424546 245854
rect 424782 245618 424866 245854
rect 425102 245618 484546 245854
rect 484782 245618 484866 245854
rect 485102 245618 544546 245854
rect 544782 245618 544866 245854
rect 545102 245618 587262 245854
rect 587498 245618 587582 245854
rect 587818 245618 588810 245854
rect -4886 245586 588810 245618
rect -2966 242454 586890 242486
rect -2966 242218 -1974 242454
rect -1738 242218 -1654 242454
rect -1418 242218 826 242454
rect 1062 242218 1146 242454
rect 1382 242218 60826 242454
rect 61062 242218 61146 242454
rect 61382 242218 120826 242454
rect 121062 242218 121146 242454
rect 121382 242218 180826 242454
rect 181062 242218 181146 242454
rect 181382 242218 204250 242454
rect 204486 242218 234970 242454
rect 235206 242218 300826 242454
rect 301062 242218 301146 242454
rect 301382 242218 360826 242454
rect 361062 242218 361146 242454
rect 361382 242218 420826 242454
rect 421062 242218 421146 242454
rect 421382 242218 480826 242454
rect 481062 242218 481146 242454
rect 481382 242218 540826 242454
rect 541062 242218 541146 242454
rect 541382 242218 585342 242454
rect 585578 242218 585662 242454
rect 585898 242218 586890 242454
rect -2966 242134 586890 242218
rect -2966 241898 -1974 242134
rect -1738 241898 -1654 242134
rect -1418 241898 826 242134
rect 1062 241898 1146 242134
rect 1382 241898 60826 242134
rect 61062 241898 61146 242134
rect 61382 241898 120826 242134
rect 121062 241898 121146 242134
rect 121382 241898 180826 242134
rect 181062 241898 181146 242134
rect 181382 241898 204250 242134
rect 204486 241898 234970 242134
rect 235206 241898 300826 242134
rect 301062 241898 301146 242134
rect 301382 241898 360826 242134
rect 361062 241898 361146 242134
rect 361382 241898 420826 242134
rect 421062 241898 421146 242134
rect 421382 241898 480826 242134
rect 481062 241898 481146 242134
rect 481382 241898 540826 242134
rect 541062 241898 541146 242134
rect 541382 241898 585342 242134
rect 585578 241898 585662 242134
rect 585898 241898 586890 242134
rect -2966 241866 586890 241898
rect -8726 223614 592650 223646
rect -8726 223378 -8694 223614
rect -8458 223378 -8374 223614
rect -8138 223378 41986 223614
rect 42222 223378 42306 223614
rect 42542 223378 101986 223614
rect 102222 223378 102306 223614
rect 102542 223378 161986 223614
rect 162222 223378 162306 223614
rect 162542 223378 281986 223614
rect 282222 223378 282306 223614
rect 282542 223378 341986 223614
rect 342222 223378 342306 223614
rect 342542 223378 401986 223614
rect 402222 223378 402306 223614
rect 402542 223378 461986 223614
rect 462222 223378 462306 223614
rect 462542 223378 521986 223614
rect 522222 223378 522306 223614
rect 522542 223378 592062 223614
rect 592298 223378 592382 223614
rect 592618 223378 592650 223614
rect -8726 223294 592650 223378
rect -8726 223058 -8694 223294
rect -8458 223058 -8374 223294
rect -8138 223058 41986 223294
rect 42222 223058 42306 223294
rect 42542 223058 101986 223294
rect 102222 223058 102306 223294
rect 102542 223058 161986 223294
rect 162222 223058 162306 223294
rect 162542 223058 281986 223294
rect 282222 223058 282306 223294
rect 282542 223058 341986 223294
rect 342222 223058 342306 223294
rect 342542 223058 401986 223294
rect 402222 223058 402306 223294
rect 402542 223058 461986 223294
rect 462222 223058 462306 223294
rect 462542 223058 521986 223294
rect 522222 223058 522306 223294
rect 522542 223058 592062 223294
rect 592298 223058 592382 223294
rect 592618 223058 592650 223294
rect -8726 223026 592650 223058
rect -6806 219894 590730 219926
rect -6806 219658 -6774 219894
rect -6538 219658 -6454 219894
rect -6218 219658 38266 219894
rect 38502 219658 38586 219894
rect 38822 219658 98266 219894
rect 98502 219658 98586 219894
rect 98822 219658 158266 219894
rect 158502 219658 158586 219894
rect 158822 219658 278266 219894
rect 278502 219658 278586 219894
rect 278822 219658 338266 219894
rect 338502 219658 338586 219894
rect 338822 219658 398266 219894
rect 398502 219658 398586 219894
rect 398822 219658 458266 219894
rect 458502 219658 458586 219894
rect 458822 219658 518266 219894
rect 518502 219658 518586 219894
rect 518822 219658 578266 219894
rect 578502 219658 578586 219894
rect 578822 219658 590142 219894
rect 590378 219658 590462 219894
rect 590698 219658 590730 219894
rect -6806 219574 590730 219658
rect -6806 219338 -6774 219574
rect -6538 219338 -6454 219574
rect -6218 219338 38266 219574
rect 38502 219338 38586 219574
rect 38822 219338 98266 219574
rect 98502 219338 98586 219574
rect 98822 219338 158266 219574
rect 158502 219338 158586 219574
rect 158822 219338 278266 219574
rect 278502 219338 278586 219574
rect 278822 219338 338266 219574
rect 338502 219338 338586 219574
rect 338822 219338 398266 219574
rect 398502 219338 398586 219574
rect 398822 219338 458266 219574
rect 458502 219338 458586 219574
rect 458822 219338 518266 219574
rect 518502 219338 518586 219574
rect 518822 219338 578266 219574
rect 578502 219338 578586 219574
rect 578822 219338 590142 219574
rect 590378 219338 590462 219574
rect 590698 219338 590730 219574
rect -6806 219306 590730 219338
rect 218156 218058 249756 218100
rect 218156 217822 218198 218058
rect 218434 217822 249478 218058
rect 249714 217822 249756 218058
rect 218156 217780 249756 217822
rect -4886 216174 588810 216206
rect -4886 215938 -4854 216174
rect -4618 215938 -4534 216174
rect -4298 215938 34546 216174
rect 34782 215938 34866 216174
rect 35102 215938 94546 216174
rect 94782 215938 94866 216174
rect 95102 215938 154546 216174
rect 154782 215938 154866 216174
rect 155102 215938 274546 216174
rect 274782 215938 274866 216174
rect 275102 215938 334546 216174
rect 334782 215938 334866 216174
rect 335102 215938 394546 216174
rect 394782 215938 394866 216174
rect 395102 215938 454546 216174
rect 454782 215938 454866 216174
rect 455102 215938 514546 216174
rect 514782 215938 514866 216174
rect 515102 215938 574546 216174
rect 574782 215938 574866 216174
rect 575102 215938 588222 216174
rect 588458 215938 588542 216174
rect 588778 215938 588810 216174
rect -4886 215854 588810 215938
rect -4886 215618 -4854 215854
rect -4618 215618 -4534 215854
rect -4298 215618 34546 215854
rect 34782 215618 34866 215854
rect 35102 215618 94546 215854
rect 94782 215618 94866 215854
rect 95102 215618 154546 215854
rect 154782 215618 154866 215854
rect 155102 215618 274546 215854
rect 274782 215618 274866 215854
rect 275102 215618 334546 215854
rect 334782 215618 334866 215854
rect 335102 215618 394546 215854
rect 394782 215618 394866 215854
rect 395102 215618 454546 215854
rect 454782 215618 454866 215854
rect 455102 215618 514546 215854
rect 514782 215618 514866 215854
rect 515102 215618 574546 215854
rect 574782 215618 574866 215854
rect 575102 215618 588222 215854
rect 588458 215618 588542 215854
rect 588778 215618 588810 215854
rect -4886 215586 588810 215618
rect -2966 212454 586890 212486
rect -2966 212218 -2934 212454
rect -2698 212218 -2614 212454
rect -2378 212218 30826 212454
rect 31062 212218 31146 212454
rect 31382 212218 90826 212454
rect 91062 212218 91146 212454
rect 91382 212218 150826 212454
rect 151062 212218 151146 212454
rect 151382 212218 219610 212454
rect 219846 212218 270826 212454
rect 271062 212218 271146 212454
rect 271382 212218 330826 212454
rect 331062 212218 331146 212454
rect 331382 212218 390826 212454
rect 391062 212218 391146 212454
rect 391382 212218 450826 212454
rect 451062 212218 451146 212454
rect 451382 212218 510826 212454
rect 511062 212218 511146 212454
rect 511382 212218 570826 212454
rect 571062 212218 571146 212454
rect 571382 212218 586302 212454
rect 586538 212218 586622 212454
rect 586858 212218 586890 212454
rect -2966 212134 586890 212218
rect -2966 211898 -2934 212134
rect -2698 211898 -2614 212134
rect -2378 211898 30826 212134
rect 31062 211898 31146 212134
rect 31382 211898 90826 212134
rect 91062 211898 91146 212134
rect 91382 211898 150826 212134
rect 151062 211898 151146 212134
rect 151382 211898 219610 212134
rect 219846 211898 270826 212134
rect 271062 211898 271146 212134
rect 271382 211898 330826 212134
rect 331062 211898 331146 212134
rect 331382 211898 390826 212134
rect 391062 211898 391146 212134
rect 391382 211898 450826 212134
rect 451062 211898 451146 212134
rect 451382 211898 510826 212134
rect 511062 211898 511146 212134
rect 511382 211898 570826 212134
rect 571062 211898 571146 212134
rect 571382 211898 586302 212134
rect 586538 211898 586622 212134
rect 586858 211898 586890 212134
rect -2966 211866 586890 211898
rect 3244 204458 249756 204500
rect 3244 204222 3286 204458
rect 3522 204222 249478 204458
rect 249714 204222 249756 204458
rect 3244 204180 249756 204222
rect -8726 193614 592650 193646
rect -8726 193378 -7734 193614
rect -7498 193378 -7414 193614
rect -7178 193378 11986 193614
rect 12222 193378 12306 193614
rect 12542 193378 71986 193614
rect 72222 193378 72306 193614
rect 72542 193378 131986 193614
rect 132222 193378 132306 193614
rect 132542 193378 191986 193614
rect 192222 193378 192306 193614
rect 192542 193378 251986 193614
rect 252222 193378 252306 193614
rect 252542 193378 311986 193614
rect 312222 193378 312306 193614
rect 312542 193378 371986 193614
rect 372222 193378 372306 193614
rect 372542 193378 431986 193614
rect 432222 193378 432306 193614
rect 432542 193378 491986 193614
rect 492222 193378 492306 193614
rect 492542 193378 551986 193614
rect 552222 193378 552306 193614
rect 552542 193378 591102 193614
rect 591338 193378 591422 193614
rect 591658 193378 592650 193614
rect -8726 193294 592650 193378
rect -8726 193058 -7734 193294
rect -7498 193058 -7414 193294
rect -7178 193058 11986 193294
rect 12222 193058 12306 193294
rect 12542 193058 71986 193294
rect 72222 193058 72306 193294
rect 72542 193058 131986 193294
rect 132222 193058 132306 193294
rect 132542 193058 191986 193294
rect 192222 193058 192306 193294
rect 192542 193058 251986 193294
rect 252222 193058 252306 193294
rect 252542 193058 311986 193294
rect 312222 193058 312306 193294
rect 312542 193058 371986 193294
rect 372222 193058 372306 193294
rect 372542 193058 431986 193294
rect 432222 193058 432306 193294
rect 432542 193058 491986 193294
rect 492222 193058 492306 193294
rect 492542 193058 551986 193294
rect 552222 193058 552306 193294
rect 552542 193058 591102 193294
rect 591338 193058 591422 193294
rect 591658 193058 592650 193294
rect -8726 193026 592650 193058
rect -6806 189894 590730 189926
rect -6806 189658 -5814 189894
rect -5578 189658 -5494 189894
rect -5258 189658 8266 189894
rect 8502 189658 8586 189894
rect 8822 189658 68266 189894
rect 68502 189658 68586 189894
rect 68822 189658 128266 189894
rect 128502 189658 128586 189894
rect 128822 189658 188266 189894
rect 188502 189658 188586 189894
rect 188822 189658 248266 189894
rect 248502 189658 248586 189894
rect 248822 189658 308266 189894
rect 308502 189658 308586 189894
rect 308822 189658 368266 189894
rect 368502 189658 368586 189894
rect 368822 189658 428266 189894
rect 428502 189658 428586 189894
rect 428822 189658 488266 189894
rect 488502 189658 488586 189894
rect 488822 189658 548266 189894
rect 548502 189658 548586 189894
rect 548822 189658 589182 189894
rect 589418 189658 589502 189894
rect 589738 189658 590730 189894
rect -6806 189574 590730 189658
rect -6806 189338 -5814 189574
rect -5578 189338 -5494 189574
rect -5258 189338 8266 189574
rect 8502 189338 8586 189574
rect 8822 189338 68266 189574
rect 68502 189338 68586 189574
rect 68822 189338 128266 189574
rect 128502 189338 128586 189574
rect 128822 189338 188266 189574
rect 188502 189338 188586 189574
rect 188822 189338 248266 189574
rect 248502 189338 248586 189574
rect 248822 189338 308266 189574
rect 308502 189338 308586 189574
rect 308822 189338 368266 189574
rect 368502 189338 368586 189574
rect 368822 189338 428266 189574
rect 428502 189338 428586 189574
rect 428822 189338 488266 189574
rect 488502 189338 488586 189574
rect 488822 189338 548266 189574
rect 548502 189338 548586 189574
rect 548822 189338 589182 189574
rect 589418 189338 589502 189574
rect 589738 189338 590730 189574
rect -6806 189306 590730 189338
rect -4886 186174 588810 186206
rect -4886 185938 -3894 186174
rect -3658 185938 -3574 186174
rect -3338 185938 4546 186174
rect 4782 185938 4866 186174
rect 5102 185938 64546 186174
rect 64782 185938 64866 186174
rect 65102 185938 124546 186174
rect 124782 185938 124866 186174
rect 125102 185938 184546 186174
rect 184782 185938 184866 186174
rect 185102 185938 244546 186174
rect 244782 185938 244866 186174
rect 245102 185938 304546 186174
rect 304782 185938 304866 186174
rect 305102 185938 364546 186174
rect 364782 185938 364866 186174
rect 365102 185938 424546 186174
rect 424782 185938 424866 186174
rect 425102 185938 484546 186174
rect 484782 185938 484866 186174
rect 485102 185938 544546 186174
rect 544782 185938 544866 186174
rect 545102 185938 587262 186174
rect 587498 185938 587582 186174
rect 587818 185938 588810 186174
rect -4886 185854 588810 185938
rect -4886 185618 -3894 185854
rect -3658 185618 -3574 185854
rect -3338 185618 4546 185854
rect 4782 185618 4866 185854
rect 5102 185618 64546 185854
rect 64782 185618 64866 185854
rect 65102 185618 124546 185854
rect 124782 185618 124866 185854
rect 125102 185618 184546 185854
rect 184782 185618 184866 185854
rect 185102 185618 244546 185854
rect 244782 185618 244866 185854
rect 245102 185618 304546 185854
rect 304782 185618 304866 185854
rect 305102 185618 364546 185854
rect 364782 185618 364866 185854
rect 365102 185618 424546 185854
rect 424782 185618 424866 185854
rect 425102 185618 484546 185854
rect 484782 185618 484866 185854
rect 485102 185618 544546 185854
rect 544782 185618 544866 185854
rect 545102 185618 587262 185854
rect 587498 185618 587582 185854
rect 587818 185618 588810 185854
rect -4886 185586 588810 185618
rect -2966 182454 586890 182486
rect -2966 182218 -1974 182454
rect -1738 182218 -1654 182454
rect -1418 182218 826 182454
rect 1062 182218 1146 182454
rect 1382 182218 60826 182454
rect 61062 182218 61146 182454
rect 61382 182218 120826 182454
rect 121062 182218 121146 182454
rect 121382 182218 180826 182454
rect 181062 182218 181146 182454
rect 181382 182218 240826 182454
rect 241062 182218 241146 182454
rect 241382 182218 300826 182454
rect 301062 182218 301146 182454
rect 301382 182218 360826 182454
rect 361062 182218 361146 182454
rect 361382 182218 420826 182454
rect 421062 182218 421146 182454
rect 421382 182218 480826 182454
rect 481062 182218 481146 182454
rect 481382 182218 540826 182454
rect 541062 182218 541146 182454
rect 541382 182218 585342 182454
rect 585578 182218 585662 182454
rect 585898 182218 586890 182454
rect -2966 182134 586890 182218
rect -2966 181898 -1974 182134
rect -1738 181898 -1654 182134
rect -1418 181898 826 182134
rect 1062 181898 1146 182134
rect 1382 181898 60826 182134
rect 61062 181898 61146 182134
rect 61382 181898 120826 182134
rect 121062 181898 121146 182134
rect 121382 181898 180826 182134
rect 181062 181898 181146 182134
rect 181382 181898 240826 182134
rect 241062 181898 241146 182134
rect 241382 181898 300826 182134
rect 301062 181898 301146 182134
rect 301382 181898 360826 182134
rect 361062 181898 361146 182134
rect 361382 181898 420826 182134
rect 421062 181898 421146 182134
rect 421382 181898 480826 182134
rect 481062 181898 481146 182134
rect 481382 181898 540826 182134
rect 541062 181898 541146 182134
rect 541382 181898 585342 182134
rect 585578 181898 585662 182134
rect 585898 181898 586890 182134
rect -2966 181866 586890 181898
rect -8726 163614 592650 163646
rect -8726 163378 -8694 163614
rect -8458 163378 -8374 163614
rect -8138 163378 41986 163614
rect 42222 163378 42306 163614
rect 42542 163378 101986 163614
rect 102222 163378 102306 163614
rect 102542 163378 161986 163614
rect 162222 163378 162306 163614
rect 162542 163378 221986 163614
rect 222222 163378 222306 163614
rect 222542 163378 281986 163614
rect 282222 163378 282306 163614
rect 282542 163378 341986 163614
rect 342222 163378 342306 163614
rect 342542 163378 401986 163614
rect 402222 163378 402306 163614
rect 402542 163378 461986 163614
rect 462222 163378 462306 163614
rect 462542 163378 521986 163614
rect 522222 163378 522306 163614
rect 522542 163378 592062 163614
rect 592298 163378 592382 163614
rect 592618 163378 592650 163614
rect -8726 163294 592650 163378
rect -8726 163058 -8694 163294
rect -8458 163058 -8374 163294
rect -8138 163058 41986 163294
rect 42222 163058 42306 163294
rect 42542 163058 101986 163294
rect 102222 163058 102306 163294
rect 102542 163058 161986 163294
rect 162222 163058 162306 163294
rect 162542 163058 221986 163294
rect 222222 163058 222306 163294
rect 222542 163058 281986 163294
rect 282222 163058 282306 163294
rect 282542 163058 341986 163294
rect 342222 163058 342306 163294
rect 342542 163058 401986 163294
rect 402222 163058 402306 163294
rect 402542 163058 461986 163294
rect 462222 163058 462306 163294
rect 462542 163058 521986 163294
rect 522222 163058 522306 163294
rect 522542 163058 592062 163294
rect 592298 163058 592382 163294
rect 592618 163058 592650 163294
rect -8726 163026 592650 163058
rect -6806 159894 590730 159926
rect -6806 159658 -6774 159894
rect -6538 159658 -6454 159894
rect -6218 159658 38266 159894
rect 38502 159658 38586 159894
rect 38822 159658 98266 159894
rect 98502 159658 98586 159894
rect 98822 159658 158266 159894
rect 158502 159658 158586 159894
rect 158822 159658 218266 159894
rect 218502 159658 218586 159894
rect 218822 159658 278266 159894
rect 278502 159658 278586 159894
rect 278822 159658 338266 159894
rect 338502 159658 338586 159894
rect 338822 159658 398266 159894
rect 398502 159658 398586 159894
rect 398822 159658 458266 159894
rect 458502 159658 458586 159894
rect 458822 159658 518266 159894
rect 518502 159658 518586 159894
rect 518822 159658 578266 159894
rect 578502 159658 578586 159894
rect 578822 159658 590142 159894
rect 590378 159658 590462 159894
rect 590698 159658 590730 159894
rect -6806 159574 590730 159658
rect -6806 159338 -6774 159574
rect -6538 159338 -6454 159574
rect -6218 159338 38266 159574
rect 38502 159338 38586 159574
rect 38822 159338 98266 159574
rect 98502 159338 98586 159574
rect 98822 159338 158266 159574
rect 158502 159338 158586 159574
rect 158822 159338 218266 159574
rect 218502 159338 218586 159574
rect 218822 159338 278266 159574
rect 278502 159338 278586 159574
rect 278822 159338 338266 159574
rect 338502 159338 338586 159574
rect 338822 159338 398266 159574
rect 398502 159338 398586 159574
rect 398822 159338 458266 159574
rect 458502 159338 458586 159574
rect 458822 159338 518266 159574
rect 518502 159338 518586 159574
rect 518822 159338 578266 159574
rect 578502 159338 578586 159574
rect 578822 159338 590142 159574
rect 590378 159338 590462 159574
rect 590698 159338 590730 159574
rect -6806 159306 590730 159338
rect -4886 156174 588810 156206
rect -4886 155938 -4854 156174
rect -4618 155938 -4534 156174
rect -4298 155938 34546 156174
rect 34782 155938 34866 156174
rect 35102 155938 94546 156174
rect 94782 155938 94866 156174
rect 95102 155938 154546 156174
rect 154782 155938 154866 156174
rect 155102 155938 214546 156174
rect 214782 155938 214866 156174
rect 215102 155938 274546 156174
rect 274782 155938 274866 156174
rect 275102 155938 334546 156174
rect 334782 155938 334866 156174
rect 335102 155938 394546 156174
rect 394782 155938 394866 156174
rect 395102 155938 454546 156174
rect 454782 155938 454866 156174
rect 455102 155938 514546 156174
rect 514782 155938 514866 156174
rect 515102 155938 574546 156174
rect 574782 155938 574866 156174
rect 575102 155938 588222 156174
rect 588458 155938 588542 156174
rect 588778 155938 588810 156174
rect -4886 155854 588810 155938
rect -4886 155618 -4854 155854
rect -4618 155618 -4534 155854
rect -4298 155618 34546 155854
rect 34782 155618 34866 155854
rect 35102 155618 94546 155854
rect 94782 155618 94866 155854
rect 95102 155618 154546 155854
rect 154782 155618 154866 155854
rect 155102 155618 214546 155854
rect 214782 155618 214866 155854
rect 215102 155618 274546 155854
rect 274782 155618 274866 155854
rect 275102 155618 334546 155854
rect 334782 155618 334866 155854
rect 335102 155618 394546 155854
rect 394782 155618 394866 155854
rect 395102 155618 454546 155854
rect 454782 155618 454866 155854
rect 455102 155618 514546 155854
rect 514782 155618 514866 155854
rect 515102 155618 574546 155854
rect 574782 155618 574866 155854
rect 575102 155618 588222 155854
rect 588458 155618 588542 155854
rect 588778 155618 588810 155854
rect -4886 155586 588810 155618
rect -2966 152454 586890 152486
rect -2966 152218 -2934 152454
rect -2698 152218 -2614 152454
rect -2378 152218 30826 152454
rect 31062 152218 31146 152454
rect 31382 152218 90826 152454
rect 91062 152218 91146 152454
rect 91382 152218 150826 152454
rect 151062 152218 151146 152454
rect 151382 152218 210826 152454
rect 211062 152218 211146 152454
rect 211382 152218 270826 152454
rect 271062 152218 271146 152454
rect 271382 152218 330826 152454
rect 331062 152218 331146 152454
rect 331382 152218 390826 152454
rect 391062 152218 391146 152454
rect 391382 152218 450826 152454
rect 451062 152218 451146 152454
rect 451382 152218 510826 152454
rect 511062 152218 511146 152454
rect 511382 152218 570826 152454
rect 571062 152218 571146 152454
rect 571382 152218 586302 152454
rect 586538 152218 586622 152454
rect 586858 152218 586890 152454
rect -2966 152134 586890 152218
rect -2966 151898 -2934 152134
rect -2698 151898 -2614 152134
rect -2378 151898 30826 152134
rect 31062 151898 31146 152134
rect 31382 151898 90826 152134
rect 91062 151898 91146 152134
rect 91382 151898 150826 152134
rect 151062 151898 151146 152134
rect 151382 151898 210826 152134
rect 211062 151898 211146 152134
rect 211382 151898 270826 152134
rect 271062 151898 271146 152134
rect 271382 151898 330826 152134
rect 331062 151898 331146 152134
rect 331382 151898 390826 152134
rect 391062 151898 391146 152134
rect 391382 151898 450826 152134
rect 451062 151898 451146 152134
rect 451382 151898 510826 152134
rect 511062 151898 511146 152134
rect 511382 151898 570826 152134
rect 571062 151898 571146 152134
rect 571382 151898 586302 152134
rect 586538 151898 586622 152134
rect 586858 151898 586890 152134
rect -2966 151866 586890 151898
rect -8726 133614 592650 133646
rect -8726 133378 -7734 133614
rect -7498 133378 -7414 133614
rect -7178 133378 11986 133614
rect 12222 133378 12306 133614
rect 12542 133378 71986 133614
rect 72222 133378 72306 133614
rect 72542 133378 131986 133614
rect 132222 133378 132306 133614
rect 132542 133378 191986 133614
rect 192222 133378 192306 133614
rect 192542 133378 251986 133614
rect 252222 133378 252306 133614
rect 252542 133378 311986 133614
rect 312222 133378 312306 133614
rect 312542 133378 371986 133614
rect 372222 133378 372306 133614
rect 372542 133378 431986 133614
rect 432222 133378 432306 133614
rect 432542 133378 491986 133614
rect 492222 133378 492306 133614
rect 492542 133378 551986 133614
rect 552222 133378 552306 133614
rect 552542 133378 591102 133614
rect 591338 133378 591422 133614
rect 591658 133378 592650 133614
rect -8726 133294 592650 133378
rect -8726 133058 -7734 133294
rect -7498 133058 -7414 133294
rect -7178 133058 11986 133294
rect 12222 133058 12306 133294
rect 12542 133058 71986 133294
rect 72222 133058 72306 133294
rect 72542 133058 131986 133294
rect 132222 133058 132306 133294
rect 132542 133058 191986 133294
rect 192222 133058 192306 133294
rect 192542 133058 251986 133294
rect 252222 133058 252306 133294
rect 252542 133058 311986 133294
rect 312222 133058 312306 133294
rect 312542 133058 371986 133294
rect 372222 133058 372306 133294
rect 372542 133058 431986 133294
rect 432222 133058 432306 133294
rect 432542 133058 491986 133294
rect 492222 133058 492306 133294
rect 492542 133058 551986 133294
rect 552222 133058 552306 133294
rect 552542 133058 591102 133294
rect 591338 133058 591422 133294
rect 591658 133058 592650 133294
rect -8726 133026 592650 133058
rect -6806 129894 590730 129926
rect -6806 129658 -5814 129894
rect -5578 129658 -5494 129894
rect -5258 129658 8266 129894
rect 8502 129658 8586 129894
rect 8822 129658 68266 129894
rect 68502 129658 68586 129894
rect 68822 129658 128266 129894
rect 128502 129658 128586 129894
rect 128822 129658 188266 129894
rect 188502 129658 188586 129894
rect 188822 129658 248266 129894
rect 248502 129658 248586 129894
rect 248822 129658 308266 129894
rect 308502 129658 308586 129894
rect 308822 129658 368266 129894
rect 368502 129658 368586 129894
rect 368822 129658 428266 129894
rect 428502 129658 428586 129894
rect 428822 129658 488266 129894
rect 488502 129658 488586 129894
rect 488822 129658 548266 129894
rect 548502 129658 548586 129894
rect 548822 129658 589182 129894
rect 589418 129658 589502 129894
rect 589738 129658 590730 129894
rect -6806 129574 590730 129658
rect -6806 129338 -5814 129574
rect -5578 129338 -5494 129574
rect -5258 129338 8266 129574
rect 8502 129338 8586 129574
rect 8822 129338 68266 129574
rect 68502 129338 68586 129574
rect 68822 129338 128266 129574
rect 128502 129338 128586 129574
rect 128822 129338 188266 129574
rect 188502 129338 188586 129574
rect 188822 129338 248266 129574
rect 248502 129338 248586 129574
rect 248822 129338 308266 129574
rect 308502 129338 308586 129574
rect 308822 129338 368266 129574
rect 368502 129338 368586 129574
rect 368822 129338 428266 129574
rect 428502 129338 428586 129574
rect 428822 129338 488266 129574
rect 488502 129338 488586 129574
rect 488822 129338 548266 129574
rect 548502 129338 548586 129574
rect 548822 129338 589182 129574
rect 589418 129338 589502 129574
rect 589738 129338 590730 129574
rect -6806 129306 590730 129338
rect -4886 126174 588810 126206
rect -4886 125938 -3894 126174
rect -3658 125938 -3574 126174
rect -3338 125938 4546 126174
rect 4782 125938 4866 126174
rect 5102 125938 64546 126174
rect 64782 125938 64866 126174
rect 65102 125938 124546 126174
rect 124782 125938 124866 126174
rect 125102 125938 184546 126174
rect 184782 125938 184866 126174
rect 185102 125938 244546 126174
rect 244782 125938 244866 126174
rect 245102 125938 304546 126174
rect 304782 125938 304866 126174
rect 305102 125938 364546 126174
rect 364782 125938 364866 126174
rect 365102 125938 424546 126174
rect 424782 125938 424866 126174
rect 425102 125938 484546 126174
rect 484782 125938 484866 126174
rect 485102 125938 544546 126174
rect 544782 125938 544866 126174
rect 545102 125938 587262 126174
rect 587498 125938 587582 126174
rect 587818 125938 588810 126174
rect -4886 125854 588810 125938
rect -4886 125618 -3894 125854
rect -3658 125618 -3574 125854
rect -3338 125618 4546 125854
rect 4782 125618 4866 125854
rect 5102 125618 64546 125854
rect 64782 125618 64866 125854
rect 65102 125618 124546 125854
rect 124782 125618 124866 125854
rect 125102 125618 184546 125854
rect 184782 125618 184866 125854
rect 185102 125618 244546 125854
rect 244782 125618 244866 125854
rect 245102 125618 304546 125854
rect 304782 125618 304866 125854
rect 305102 125618 364546 125854
rect 364782 125618 364866 125854
rect 365102 125618 424546 125854
rect 424782 125618 424866 125854
rect 425102 125618 484546 125854
rect 484782 125618 484866 125854
rect 485102 125618 544546 125854
rect 544782 125618 544866 125854
rect 545102 125618 587262 125854
rect 587498 125618 587582 125854
rect 587818 125618 588810 125854
rect -4886 125586 588810 125618
rect -2966 122454 586890 122486
rect -2966 122218 -1974 122454
rect -1738 122218 -1654 122454
rect -1418 122218 826 122454
rect 1062 122218 1146 122454
rect 1382 122218 60826 122454
rect 61062 122218 61146 122454
rect 61382 122218 120826 122454
rect 121062 122218 121146 122454
rect 121382 122218 180826 122454
rect 181062 122218 181146 122454
rect 181382 122218 240826 122454
rect 241062 122218 241146 122454
rect 241382 122218 300826 122454
rect 301062 122218 301146 122454
rect 301382 122218 360826 122454
rect 361062 122218 361146 122454
rect 361382 122218 420826 122454
rect 421062 122218 421146 122454
rect 421382 122218 480826 122454
rect 481062 122218 481146 122454
rect 481382 122218 540826 122454
rect 541062 122218 541146 122454
rect 541382 122218 585342 122454
rect 585578 122218 585662 122454
rect 585898 122218 586890 122454
rect -2966 122134 586890 122218
rect -2966 121898 -1974 122134
rect -1738 121898 -1654 122134
rect -1418 121898 826 122134
rect 1062 121898 1146 122134
rect 1382 121898 60826 122134
rect 61062 121898 61146 122134
rect 61382 121898 120826 122134
rect 121062 121898 121146 122134
rect 121382 121898 180826 122134
rect 181062 121898 181146 122134
rect 181382 121898 240826 122134
rect 241062 121898 241146 122134
rect 241382 121898 300826 122134
rect 301062 121898 301146 122134
rect 301382 121898 360826 122134
rect 361062 121898 361146 122134
rect 361382 121898 420826 122134
rect 421062 121898 421146 122134
rect 421382 121898 480826 122134
rect 481062 121898 481146 122134
rect 481382 121898 540826 122134
rect 541062 121898 541146 122134
rect 541382 121898 585342 122134
rect 585578 121898 585662 122134
rect 585898 121898 586890 122134
rect -2966 121866 586890 121898
rect -8726 103614 592650 103646
rect -8726 103378 -8694 103614
rect -8458 103378 -8374 103614
rect -8138 103378 41986 103614
rect 42222 103378 42306 103614
rect 42542 103378 101986 103614
rect 102222 103378 102306 103614
rect 102542 103378 161986 103614
rect 162222 103378 162306 103614
rect 162542 103378 221986 103614
rect 222222 103378 222306 103614
rect 222542 103378 281986 103614
rect 282222 103378 282306 103614
rect 282542 103378 341986 103614
rect 342222 103378 342306 103614
rect 342542 103378 401986 103614
rect 402222 103378 402306 103614
rect 402542 103378 461986 103614
rect 462222 103378 462306 103614
rect 462542 103378 521986 103614
rect 522222 103378 522306 103614
rect 522542 103378 592062 103614
rect 592298 103378 592382 103614
rect 592618 103378 592650 103614
rect -8726 103294 592650 103378
rect -8726 103058 -8694 103294
rect -8458 103058 -8374 103294
rect -8138 103058 41986 103294
rect 42222 103058 42306 103294
rect 42542 103058 101986 103294
rect 102222 103058 102306 103294
rect 102542 103058 161986 103294
rect 162222 103058 162306 103294
rect 162542 103058 221986 103294
rect 222222 103058 222306 103294
rect 222542 103058 281986 103294
rect 282222 103058 282306 103294
rect 282542 103058 341986 103294
rect 342222 103058 342306 103294
rect 342542 103058 401986 103294
rect 402222 103058 402306 103294
rect 402542 103058 461986 103294
rect 462222 103058 462306 103294
rect 462542 103058 521986 103294
rect 522222 103058 522306 103294
rect 522542 103058 592062 103294
rect 592298 103058 592382 103294
rect 592618 103058 592650 103294
rect -8726 103026 592650 103058
rect -6806 99894 590730 99926
rect -6806 99658 -6774 99894
rect -6538 99658 -6454 99894
rect -6218 99658 38266 99894
rect 38502 99658 38586 99894
rect 38822 99658 98266 99894
rect 98502 99658 98586 99894
rect 98822 99658 158266 99894
rect 158502 99658 158586 99894
rect 158822 99658 218266 99894
rect 218502 99658 218586 99894
rect 218822 99658 278266 99894
rect 278502 99658 278586 99894
rect 278822 99658 338266 99894
rect 338502 99658 338586 99894
rect 338822 99658 398266 99894
rect 398502 99658 398586 99894
rect 398822 99658 458266 99894
rect 458502 99658 458586 99894
rect 458822 99658 518266 99894
rect 518502 99658 518586 99894
rect 518822 99658 578266 99894
rect 578502 99658 578586 99894
rect 578822 99658 590142 99894
rect 590378 99658 590462 99894
rect 590698 99658 590730 99894
rect -6806 99574 590730 99658
rect -6806 99338 -6774 99574
rect -6538 99338 -6454 99574
rect -6218 99338 38266 99574
rect 38502 99338 38586 99574
rect 38822 99338 98266 99574
rect 98502 99338 98586 99574
rect 98822 99338 158266 99574
rect 158502 99338 158586 99574
rect 158822 99338 218266 99574
rect 218502 99338 218586 99574
rect 218822 99338 278266 99574
rect 278502 99338 278586 99574
rect 278822 99338 338266 99574
rect 338502 99338 338586 99574
rect 338822 99338 398266 99574
rect 398502 99338 398586 99574
rect 398822 99338 458266 99574
rect 458502 99338 458586 99574
rect 458822 99338 518266 99574
rect 518502 99338 518586 99574
rect 518822 99338 578266 99574
rect 578502 99338 578586 99574
rect 578822 99338 590142 99574
rect 590378 99338 590462 99574
rect 590698 99338 590730 99574
rect -6806 99306 590730 99338
rect -4886 96174 588810 96206
rect -4886 95938 -4854 96174
rect -4618 95938 -4534 96174
rect -4298 95938 34546 96174
rect 34782 95938 34866 96174
rect 35102 95938 94546 96174
rect 94782 95938 94866 96174
rect 95102 95938 154546 96174
rect 154782 95938 154866 96174
rect 155102 95938 214546 96174
rect 214782 95938 214866 96174
rect 215102 95938 274546 96174
rect 274782 95938 274866 96174
rect 275102 95938 334546 96174
rect 334782 95938 334866 96174
rect 335102 95938 394546 96174
rect 394782 95938 394866 96174
rect 395102 95938 454546 96174
rect 454782 95938 454866 96174
rect 455102 95938 514546 96174
rect 514782 95938 514866 96174
rect 515102 95938 574546 96174
rect 574782 95938 574866 96174
rect 575102 95938 588222 96174
rect 588458 95938 588542 96174
rect 588778 95938 588810 96174
rect -4886 95854 588810 95938
rect -4886 95618 -4854 95854
rect -4618 95618 -4534 95854
rect -4298 95618 34546 95854
rect 34782 95618 34866 95854
rect 35102 95618 94546 95854
rect 94782 95618 94866 95854
rect 95102 95618 154546 95854
rect 154782 95618 154866 95854
rect 155102 95618 214546 95854
rect 214782 95618 214866 95854
rect 215102 95618 274546 95854
rect 274782 95618 274866 95854
rect 275102 95618 334546 95854
rect 334782 95618 334866 95854
rect 335102 95618 394546 95854
rect 394782 95618 394866 95854
rect 395102 95618 454546 95854
rect 454782 95618 454866 95854
rect 455102 95618 514546 95854
rect 514782 95618 514866 95854
rect 515102 95618 574546 95854
rect 574782 95618 574866 95854
rect 575102 95618 588222 95854
rect 588458 95618 588542 95854
rect 588778 95618 588810 95854
rect -4886 95586 588810 95618
rect -2966 92454 586890 92486
rect -2966 92218 -2934 92454
rect -2698 92218 -2614 92454
rect -2378 92218 30826 92454
rect 31062 92218 31146 92454
rect 31382 92218 90826 92454
rect 91062 92218 91146 92454
rect 91382 92218 150826 92454
rect 151062 92218 151146 92454
rect 151382 92218 210826 92454
rect 211062 92218 211146 92454
rect 211382 92218 270826 92454
rect 271062 92218 271146 92454
rect 271382 92218 330826 92454
rect 331062 92218 331146 92454
rect 331382 92218 390826 92454
rect 391062 92218 391146 92454
rect 391382 92218 450826 92454
rect 451062 92218 451146 92454
rect 451382 92218 510826 92454
rect 511062 92218 511146 92454
rect 511382 92218 570826 92454
rect 571062 92218 571146 92454
rect 571382 92218 586302 92454
rect 586538 92218 586622 92454
rect 586858 92218 586890 92454
rect -2966 92134 586890 92218
rect -2966 91898 -2934 92134
rect -2698 91898 -2614 92134
rect -2378 91898 30826 92134
rect 31062 91898 31146 92134
rect 31382 91898 90826 92134
rect 91062 91898 91146 92134
rect 91382 91898 150826 92134
rect 151062 91898 151146 92134
rect 151382 91898 210826 92134
rect 211062 91898 211146 92134
rect 211382 91898 270826 92134
rect 271062 91898 271146 92134
rect 271382 91898 330826 92134
rect 331062 91898 331146 92134
rect 331382 91898 390826 92134
rect 391062 91898 391146 92134
rect 391382 91898 450826 92134
rect 451062 91898 451146 92134
rect 451382 91898 510826 92134
rect 511062 91898 511146 92134
rect 511382 91898 570826 92134
rect 571062 91898 571146 92134
rect 571382 91898 586302 92134
rect 586538 91898 586622 92134
rect 586858 91898 586890 92134
rect -2966 91866 586890 91898
rect -8726 73614 592650 73646
rect -8726 73378 -7734 73614
rect -7498 73378 -7414 73614
rect -7178 73378 11986 73614
rect 12222 73378 12306 73614
rect 12542 73378 71986 73614
rect 72222 73378 72306 73614
rect 72542 73378 131986 73614
rect 132222 73378 132306 73614
rect 132542 73378 191986 73614
rect 192222 73378 192306 73614
rect 192542 73378 251986 73614
rect 252222 73378 252306 73614
rect 252542 73378 311986 73614
rect 312222 73378 312306 73614
rect 312542 73378 371986 73614
rect 372222 73378 372306 73614
rect 372542 73378 431986 73614
rect 432222 73378 432306 73614
rect 432542 73378 491986 73614
rect 492222 73378 492306 73614
rect 492542 73378 551986 73614
rect 552222 73378 552306 73614
rect 552542 73378 591102 73614
rect 591338 73378 591422 73614
rect 591658 73378 592650 73614
rect -8726 73294 592650 73378
rect -8726 73058 -7734 73294
rect -7498 73058 -7414 73294
rect -7178 73058 11986 73294
rect 12222 73058 12306 73294
rect 12542 73058 71986 73294
rect 72222 73058 72306 73294
rect 72542 73058 131986 73294
rect 132222 73058 132306 73294
rect 132542 73058 191986 73294
rect 192222 73058 192306 73294
rect 192542 73058 251986 73294
rect 252222 73058 252306 73294
rect 252542 73058 311986 73294
rect 312222 73058 312306 73294
rect 312542 73058 371986 73294
rect 372222 73058 372306 73294
rect 372542 73058 431986 73294
rect 432222 73058 432306 73294
rect 432542 73058 491986 73294
rect 492222 73058 492306 73294
rect 492542 73058 551986 73294
rect 552222 73058 552306 73294
rect 552542 73058 591102 73294
rect 591338 73058 591422 73294
rect 591658 73058 592650 73294
rect -8726 73026 592650 73058
rect -6806 69894 590730 69926
rect -6806 69658 -5814 69894
rect -5578 69658 -5494 69894
rect -5258 69658 8266 69894
rect 8502 69658 8586 69894
rect 8822 69658 68266 69894
rect 68502 69658 68586 69894
rect 68822 69658 128266 69894
rect 128502 69658 128586 69894
rect 128822 69658 188266 69894
rect 188502 69658 188586 69894
rect 188822 69658 248266 69894
rect 248502 69658 248586 69894
rect 248822 69658 308266 69894
rect 308502 69658 308586 69894
rect 308822 69658 368266 69894
rect 368502 69658 368586 69894
rect 368822 69658 428266 69894
rect 428502 69658 428586 69894
rect 428822 69658 488266 69894
rect 488502 69658 488586 69894
rect 488822 69658 548266 69894
rect 548502 69658 548586 69894
rect 548822 69658 589182 69894
rect 589418 69658 589502 69894
rect 589738 69658 590730 69894
rect -6806 69574 590730 69658
rect -6806 69338 -5814 69574
rect -5578 69338 -5494 69574
rect -5258 69338 8266 69574
rect 8502 69338 8586 69574
rect 8822 69338 68266 69574
rect 68502 69338 68586 69574
rect 68822 69338 128266 69574
rect 128502 69338 128586 69574
rect 128822 69338 188266 69574
rect 188502 69338 188586 69574
rect 188822 69338 248266 69574
rect 248502 69338 248586 69574
rect 248822 69338 308266 69574
rect 308502 69338 308586 69574
rect 308822 69338 368266 69574
rect 368502 69338 368586 69574
rect 368822 69338 428266 69574
rect 428502 69338 428586 69574
rect 428822 69338 488266 69574
rect 488502 69338 488586 69574
rect 488822 69338 548266 69574
rect 548502 69338 548586 69574
rect 548822 69338 589182 69574
rect 589418 69338 589502 69574
rect 589738 69338 590730 69574
rect -6806 69306 590730 69338
rect -4886 66174 588810 66206
rect -4886 65938 -3894 66174
rect -3658 65938 -3574 66174
rect -3338 65938 4546 66174
rect 4782 65938 4866 66174
rect 5102 65938 64546 66174
rect 64782 65938 64866 66174
rect 65102 65938 124546 66174
rect 124782 65938 124866 66174
rect 125102 65938 184546 66174
rect 184782 65938 184866 66174
rect 185102 65938 244546 66174
rect 244782 65938 244866 66174
rect 245102 65938 304546 66174
rect 304782 65938 304866 66174
rect 305102 65938 364546 66174
rect 364782 65938 364866 66174
rect 365102 65938 424546 66174
rect 424782 65938 424866 66174
rect 425102 65938 484546 66174
rect 484782 65938 484866 66174
rect 485102 65938 544546 66174
rect 544782 65938 544866 66174
rect 545102 65938 587262 66174
rect 587498 65938 587582 66174
rect 587818 65938 588810 66174
rect -4886 65854 588810 65938
rect -4886 65618 -3894 65854
rect -3658 65618 -3574 65854
rect -3338 65618 4546 65854
rect 4782 65618 4866 65854
rect 5102 65618 64546 65854
rect 64782 65618 64866 65854
rect 65102 65618 124546 65854
rect 124782 65618 124866 65854
rect 125102 65618 184546 65854
rect 184782 65618 184866 65854
rect 185102 65618 244546 65854
rect 244782 65618 244866 65854
rect 245102 65618 304546 65854
rect 304782 65618 304866 65854
rect 305102 65618 364546 65854
rect 364782 65618 364866 65854
rect 365102 65618 424546 65854
rect 424782 65618 424866 65854
rect 425102 65618 484546 65854
rect 484782 65618 484866 65854
rect 485102 65618 544546 65854
rect 544782 65618 544866 65854
rect 545102 65618 587262 65854
rect 587498 65618 587582 65854
rect 587818 65618 588810 65854
rect -4886 65586 588810 65618
rect -2966 62454 586890 62486
rect -2966 62218 -1974 62454
rect -1738 62218 -1654 62454
rect -1418 62218 826 62454
rect 1062 62218 1146 62454
rect 1382 62218 60826 62454
rect 61062 62218 61146 62454
rect 61382 62218 120826 62454
rect 121062 62218 121146 62454
rect 121382 62218 180826 62454
rect 181062 62218 181146 62454
rect 181382 62218 240826 62454
rect 241062 62218 241146 62454
rect 241382 62218 300826 62454
rect 301062 62218 301146 62454
rect 301382 62218 360826 62454
rect 361062 62218 361146 62454
rect 361382 62218 420826 62454
rect 421062 62218 421146 62454
rect 421382 62218 480826 62454
rect 481062 62218 481146 62454
rect 481382 62218 540826 62454
rect 541062 62218 541146 62454
rect 541382 62218 585342 62454
rect 585578 62218 585662 62454
rect 585898 62218 586890 62454
rect -2966 62134 586890 62218
rect -2966 61898 -1974 62134
rect -1738 61898 -1654 62134
rect -1418 61898 826 62134
rect 1062 61898 1146 62134
rect 1382 61898 60826 62134
rect 61062 61898 61146 62134
rect 61382 61898 120826 62134
rect 121062 61898 121146 62134
rect 121382 61898 180826 62134
rect 181062 61898 181146 62134
rect 181382 61898 240826 62134
rect 241062 61898 241146 62134
rect 241382 61898 300826 62134
rect 301062 61898 301146 62134
rect 301382 61898 360826 62134
rect 361062 61898 361146 62134
rect 361382 61898 420826 62134
rect 421062 61898 421146 62134
rect 421382 61898 480826 62134
rect 481062 61898 481146 62134
rect 481382 61898 540826 62134
rect 541062 61898 541146 62134
rect 541382 61898 585342 62134
rect 585578 61898 585662 62134
rect 585898 61898 586890 62134
rect -2966 61866 586890 61898
rect -8726 43614 592650 43646
rect -8726 43378 -8694 43614
rect -8458 43378 -8374 43614
rect -8138 43378 41986 43614
rect 42222 43378 42306 43614
rect 42542 43378 101986 43614
rect 102222 43378 102306 43614
rect 102542 43378 161986 43614
rect 162222 43378 162306 43614
rect 162542 43378 221986 43614
rect 222222 43378 222306 43614
rect 222542 43378 281986 43614
rect 282222 43378 282306 43614
rect 282542 43378 341986 43614
rect 342222 43378 342306 43614
rect 342542 43378 401986 43614
rect 402222 43378 402306 43614
rect 402542 43378 461986 43614
rect 462222 43378 462306 43614
rect 462542 43378 521986 43614
rect 522222 43378 522306 43614
rect 522542 43378 592062 43614
rect 592298 43378 592382 43614
rect 592618 43378 592650 43614
rect -8726 43294 592650 43378
rect -8726 43058 -8694 43294
rect -8458 43058 -8374 43294
rect -8138 43058 41986 43294
rect 42222 43058 42306 43294
rect 42542 43058 101986 43294
rect 102222 43058 102306 43294
rect 102542 43058 161986 43294
rect 162222 43058 162306 43294
rect 162542 43058 221986 43294
rect 222222 43058 222306 43294
rect 222542 43058 281986 43294
rect 282222 43058 282306 43294
rect 282542 43058 341986 43294
rect 342222 43058 342306 43294
rect 342542 43058 401986 43294
rect 402222 43058 402306 43294
rect 402542 43058 461986 43294
rect 462222 43058 462306 43294
rect 462542 43058 521986 43294
rect 522222 43058 522306 43294
rect 522542 43058 592062 43294
rect 592298 43058 592382 43294
rect 592618 43058 592650 43294
rect -8726 43026 592650 43058
rect -6806 39894 590730 39926
rect -6806 39658 -6774 39894
rect -6538 39658 -6454 39894
rect -6218 39658 38266 39894
rect 38502 39658 38586 39894
rect 38822 39658 98266 39894
rect 98502 39658 98586 39894
rect 98822 39658 158266 39894
rect 158502 39658 158586 39894
rect 158822 39658 218266 39894
rect 218502 39658 218586 39894
rect 218822 39658 278266 39894
rect 278502 39658 278586 39894
rect 278822 39658 338266 39894
rect 338502 39658 338586 39894
rect 338822 39658 398266 39894
rect 398502 39658 398586 39894
rect 398822 39658 458266 39894
rect 458502 39658 458586 39894
rect 458822 39658 518266 39894
rect 518502 39658 518586 39894
rect 518822 39658 578266 39894
rect 578502 39658 578586 39894
rect 578822 39658 590142 39894
rect 590378 39658 590462 39894
rect 590698 39658 590730 39894
rect -6806 39574 590730 39658
rect -6806 39338 -6774 39574
rect -6538 39338 -6454 39574
rect -6218 39338 38266 39574
rect 38502 39338 38586 39574
rect 38822 39338 98266 39574
rect 98502 39338 98586 39574
rect 98822 39338 158266 39574
rect 158502 39338 158586 39574
rect 158822 39338 218266 39574
rect 218502 39338 218586 39574
rect 218822 39338 278266 39574
rect 278502 39338 278586 39574
rect 278822 39338 338266 39574
rect 338502 39338 338586 39574
rect 338822 39338 398266 39574
rect 398502 39338 398586 39574
rect 398822 39338 458266 39574
rect 458502 39338 458586 39574
rect 458822 39338 518266 39574
rect 518502 39338 518586 39574
rect 518822 39338 578266 39574
rect 578502 39338 578586 39574
rect 578822 39338 590142 39574
rect 590378 39338 590462 39574
rect 590698 39338 590730 39574
rect -6806 39306 590730 39338
rect -4886 36174 588810 36206
rect -4886 35938 -4854 36174
rect -4618 35938 -4534 36174
rect -4298 35938 34546 36174
rect 34782 35938 34866 36174
rect 35102 35938 94546 36174
rect 94782 35938 94866 36174
rect 95102 35938 154546 36174
rect 154782 35938 154866 36174
rect 155102 35938 214546 36174
rect 214782 35938 214866 36174
rect 215102 35938 274546 36174
rect 274782 35938 274866 36174
rect 275102 35938 334546 36174
rect 334782 35938 334866 36174
rect 335102 35938 394546 36174
rect 394782 35938 394866 36174
rect 395102 35938 454546 36174
rect 454782 35938 454866 36174
rect 455102 35938 514546 36174
rect 514782 35938 514866 36174
rect 515102 35938 574546 36174
rect 574782 35938 574866 36174
rect 575102 35938 588222 36174
rect 588458 35938 588542 36174
rect 588778 35938 588810 36174
rect -4886 35854 588810 35938
rect -4886 35618 -4854 35854
rect -4618 35618 -4534 35854
rect -4298 35618 34546 35854
rect 34782 35618 34866 35854
rect 35102 35618 94546 35854
rect 94782 35618 94866 35854
rect 95102 35618 154546 35854
rect 154782 35618 154866 35854
rect 155102 35618 214546 35854
rect 214782 35618 214866 35854
rect 215102 35618 274546 35854
rect 274782 35618 274866 35854
rect 275102 35618 334546 35854
rect 334782 35618 334866 35854
rect 335102 35618 394546 35854
rect 394782 35618 394866 35854
rect 395102 35618 454546 35854
rect 454782 35618 454866 35854
rect 455102 35618 514546 35854
rect 514782 35618 514866 35854
rect 515102 35618 574546 35854
rect 574782 35618 574866 35854
rect 575102 35618 588222 35854
rect 588458 35618 588542 35854
rect 588778 35618 588810 35854
rect -4886 35586 588810 35618
rect -2966 32454 586890 32486
rect -2966 32218 -2934 32454
rect -2698 32218 -2614 32454
rect -2378 32218 30826 32454
rect 31062 32218 31146 32454
rect 31382 32218 90826 32454
rect 91062 32218 91146 32454
rect 91382 32218 150826 32454
rect 151062 32218 151146 32454
rect 151382 32218 210826 32454
rect 211062 32218 211146 32454
rect 211382 32218 270826 32454
rect 271062 32218 271146 32454
rect 271382 32218 330826 32454
rect 331062 32218 331146 32454
rect 331382 32218 390826 32454
rect 391062 32218 391146 32454
rect 391382 32218 450826 32454
rect 451062 32218 451146 32454
rect 451382 32218 510826 32454
rect 511062 32218 511146 32454
rect 511382 32218 570826 32454
rect 571062 32218 571146 32454
rect 571382 32218 586302 32454
rect 586538 32218 586622 32454
rect 586858 32218 586890 32454
rect -2966 32134 586890 32218
rect -2966 31898 -2934 32134
rect -2698 31898 -2614 32134
rect -2378 31898 30826 32134
rect 31062 31898 31146 32134
rect 31382 31898 90826 32134
rect 91062 31898 91146 32134
rect 91382 31898 150826 32134
rect 151062 31898 151146 32134
rect 151382 31898 210826 32134
rect 211062 31898 211146 32134
rect 211382 31898 270826 32134
rect 271062 31898 271146 32134
rect 271382 31898 330826 32134
rect 331062 31898 331146 32134
rect 331382 31898 390826 32134
rect 391062 31898 391146 32134
rect 391382 31898 450826 32134
rect 451062 31898 451146 32134
rect 451382 31898 510826 32134
rect 511062 31898 511146 32134
rect 511382 31898 570826 32134
rect 571062 31898 571146 32134
rect 571382 31898 586302 32134
rect 586538 31898 586622 32134
rect 586858 31898 586890 32134
rect -2966 31866 586890 31898
rect -8726 13614 592650 13646
rect -8726 13378 -7734 13614
rect -7498 13378 -7414 13614
rect -7178 13378 11986 13614
rect 12222 13378 12306 13614
rect 12542 13378 71986 13614
rect 72222 13378 72306 13614
rect 72542 13378 131986 13614
rect 132222 13378 132306 13614
rect 132542 13378 191986 13614
rect 192222 13378 192306 13614
rect 192542 13378 251986 13614
rect 252222 13378 252306 13614
rect 252542 13378 311986 13614
rect 312222 13378 312306 13614
rect 312542 13378 371986 13614
rect 372222 13378 372306 13614
rect 372542 13378 431986 13614
rect 432222 13378 432306 13614
rect 432542 13378 491986 13614
rect 492222 13378 492306 13614
rect 492542 13378 551986 13614
rect 552222 13378 552306 13614
rect 552542 13378 591102 13614
rect 591338 13378 591422 13614
rect 591658 13378 592650 13614
rect -8726 13294 592650 13378
rect -8726 13058 -7734 13294
rect -7498 13058 -7414 13294
rect -7178 13058 11986 13294
rect 12222 13058 12306 13294
rect 12542 13058 71986 13294
rect 72222 13058 72306 13294
rect 72542 13058 131986 13294
rect 132222 13058 132306 13294
rect 132542 13058 191986 13294
rect 192222 13058 192306 13294
rect 192542 13058 251986 13294
rect 252222 13058 252306 13294
rect 252542 13058 311986 13294
rect 312222 13058 312306 13294
rect 312542 13058 371986 13294
rect 372222 13058 372306 13294
rect 372542 13058 431986 13294
rect 432222 13058 432306 13294
rect 432542 13058 491986 13294
rect 492222 13058 492306 13294
rect 492542 13058 551986 13294
rect 552222 13058 552306 13294
rect 552542 13058 591102 13294
rect 591338 13058 591422 13294
rect 591658 13058 592650 13294
rect -8726 13026 592650 13058
rect -6806 9894 590730 9926
rect -6806 9658 -5814 9894
rect -5578 9658 -5494 9894
rect -5258 9658 8266 9894
rect 8502 9658 8586 9894
rect 8822 9658 68266 9894
rect 68502 9658 68586 9894
rect 68822 9658 128266 9894
rect 128502 9658 128586 9894
rect 128822 9658 188266 9894
rect 188502 9658 188586 9894
rect 188822 9658 248266 9894
rect 248502 9658 248586 9894
rect 248822 9658 308266 9894
rect 308502 9658 308586 9894
rect 308822 9658 368266 9894
rect 368502 9658 368586 9894
rect 368822 9658 428266 9894
rect 428502 9658 428586 9894
rect 428822 9658 488266 9894
rect 488502 9658 488586 9894
rect 488822 9658 548266 9894
rect 548502 9658 548586 9894
rect 548822 9658 589182 9894
rect 589418 9658 589502 9894
rect 589738 9658 590730 9894
rect -6806 9574 590730 9658
rect -6806 9338 -5814 9574
rect -5578 9338 -5494 9574
rect -5258 9338 8266 9574
rect 8502 9338 8586 9574
rect 8822 9338 68266 9574
rect 68502 9338 68586 9574
rect 68822 9338 128266 9574
rect 128502 9338 128586 9574
rect 128822 9338 188266 9574
rect 188502 9338 188586 9574
rect 188822 9338 248266 9574
rect 248502 9338 248586 9574
rect 248822 9338 308266 9574
rect 308502 9338 308586 9574
rect 308822 9338 368266 9574
rect 368502 9338 368586 9574
rect 368822 9338 428266 9574
rect 428502 9338 428586 9574
rect 428822 9338 488266 9574
rect 488502 9338 488586 9574
rect 488822 9338 548266 9574
rect 548502 9338 548586 9574
rect 548822 9338 589182 9574
rect 589418 9338 589502 9574
rect 589738 9338 590730 9574
rect -6806 9306 590730 9338
rect -4886 6174 588810 6206
rect -4886 5938 -3894 6174
rect -3658 5938 -3574 6174
rect -3338 5938 4546 6174
rect 4782 5938 4866 6174
rect 5102 5938 64546 6174
rect 64782 5938 64866 6174
rect 65102 5938 124546 6174
rect 124782 5938 124866 6174
rect 125102 5938 184546 6174
rect 184782 5938 184866 6174
rect 185102 5938 244546 6174
rect 244782 5938 244866 6174
rect 245102 5938 304546 6174
rect 304782 5938 304866 6174
rect 305102 5938 364546 6174
rect 364782 5938 364866 6174
rect 365102 5938 424546 6174
rect 424782 5938 424866 6174
rect 425102 5938 484546 6174
rect 484782 5938 484866 6174
rect 485102 5938 544546 6174
rect 544782 5938 544866 6174
rect 545102 5938 587262 6174
rect 587498 5938 587582 6174
rect 587818 5938 588810 6174
rect -4886 5854 588810 5938
rect -4886 5618 -3894 5854
rect -3658 5618 -3574 5854
rect -3338 5618 4546 5854
rect 4782 5618 4866 5854
rect 5102 5618 64546 5854
rect 64782 5618 64866 5854
rect 65102 5618 124546 5854
rect 124782 5618 124866 5854
rect 125102 5618 184546 5854
rect 184782 5618 184866 5854
rect 185102 5618 244546 5854
rect 244782 5618 244866 5854
rect 245102 5618 304546 5854
rect 304782 5618 304866 5854
rect 305102 5618 364546 5854
rect 364782 5618 364866 5854
rect 365102 5618 424546 5854
rect 424782 5618 424866 5854
rect 425102 5618 484546 5854
rect 484782 5618 484866 5854
rect 485102 5618 544546 5854
rect 544782 5618 544866 5854
rect 545102 5618 587262 5854
rect 587498 5618 587582 5854
rect 587818 5618 588810 5854
rect -4886 5586 588810 5618
rect -2966 2454 586890 2486
rect -2966 2218 -1974 2454
rect -1738 2218 -1654 2454
rect -1418 2218 826 2454
rect 1062 2218 1146 2454
rect 1382 2218 60826 2454
rect 61062 2218 61146 2454
rect 61382 2218 120826 2454
rect 121062 2218 121146 2454
rect 121382 2218 180826 2454
rect 181062 2218 181146 2454
rect 181382 2218 240826 2454
rect 241062 2218 241146 2454
rect 241382 2218 300826 2454
rect 301062 2218 301146 2454
rect 301382 2218 360826 2454
rect 361062 2218 361146 2454
rect 361382 2218 420826 2454
rect 421062 2218 421146 2454
rect 421382 2218 480826 2454
rect 481062 2218 481146 2454
rect 481382 2218 540826 2454
rect 541062 2218 541146 2454
rect 541382 2218 585342 2454
rect 585578 2218 585662 2454
rect 585898 2218 586890 2454
rect -2966 2134 586890 2218
rect -2966 1898 -1974 2134
rect -1738 1898 -1654 2134
rect -1418 1898 826 2134
rect 1062 1898 1146 2134
rect 1382 1898 60826 2134
rect 61062 1898 61146 2134
rect 61382 1898 120826 2134
rect 121062 1898 121146 2134
rect 121382 1898 180826 2134
rect 181062 1898 181146 2134
rect 181382 1898 240826 2134
rect 241062 1898 241146 2134
rect 241382 1898 300826 2134
rect 301062 1898 301146 2134
rect 301382 1898 360826 2134
rect 361062 1898 361146 2134
rect 361382 1898 420826 2134
rect 421062 1898 421146 2134
rect 421382 1898 480826 2134
rect 481062 1898 481146 2134
rect 481382 1898 540826 2134
rect 541062 1898 541146 2134
rect 541382 1898 585342 2134
rect 585578 1898 585662 2134
rect 585898 1898 586890 2134
rect -2966 1866 586890 1898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 826 -346
rect 1062 -582 1146 -346
rect 1382 -582 60826 -346
rect 61062 -582 61146 -346
rect 61382 -582 120826 -346
rect 121062 -582 121146 -346
rect 121382 -582 180826 -346
rect 181062 -582 181146 -346
rect 181382 -582 240826 -346
rect 241062 -582 241146 -346
rect 241382 -582 300826 -346
rect 301062 -582 301146 -346
rect 301382 -582 360826 -346
rect 361062 -582 361146 -346
rect 361382 -582 420826 -346
rect 421062 -582 421146 -346
rect 421382 -582 480826 -346
rect 481062 -582 481146 -346
rect 481382 -582 540826 -346
rect 541062 -582 541146 -346
rect 541382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 826 -666
rect 1062 -902 1146 -666
rect 1382 -902 60826 -666
rect 61062 -902 61146 -666
rect 61382 -902 120826 -666
rect 121062 -902 121146 -666
rect 121382 -902 180826 -666
rect 181062 -902 181146 -666
rect 181382 -902 240826 -666
rect 241062 -902 241146 -666
rect 241382 -902 300826 -666
rect 301062 -902 301146 -666
rect 301382 -902 360826 -666
rect 361062 -902 361146 -666
rect 361382 -902 420826 -666
rect 421062 -902 421146 -666
rect 421382 -902 480826 -666
rect 481062 -902 481146 -666
rect 481382 -902 540826 -666
rect 541062 -902 541146 -666
rect 541382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 30826 -1306
rect 31062 -1542 31146 -1306
rect 31382 -1542 90826 -1306
rect 91062 -1542 91146 -1306
rect 91382 -1542 150826 -1306
rect 151062 -1542 151146 -1306
rect 151382 -1542 210826 -1306
rect 211062 -1542 211146 -1306
rect 211382 -1542 270826 -1306
rect 271062 -1542 271146 -1306
rect 271382 -1542 330826 -1306
rect 331062 -1542 331146 -1306
rect 331382 -1542 390826 -1306
rect 391062 -1542 391146 -1306
rect 391382 -1542 450826 -1306
rect 451062 -1542 451146 -1306
rect 451382 -1542 510826 -1306
rect 511062 -1542 511146 -1306
rect 511382 -1542 570826 -1306
rect 571062 -1542 571146 -1306
rect 571382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 30826 -1626
rect 31062 -1862 31146 -1626
rect 31382 -1862 90826 -1626
rect 91062 -1862 91146 -1626
rect 91382 -1862 150826 -1626
rect 151062 -1862 151146 -1626
rect 151382 -1862 210826 -1626
rect 211062 -1862 211146 -1626
rect 211382 -1862 270826 -1626
rect 271062 -1862 271146 -1626
rect 271382 -1862 330826 -1626
rect 331062 -1862 331146 -1626
rect 331382 -1862 390826 -1626
rect 391062 -1862 391146 -1626
rect 391382 -1862 450826 -1626
rect 451062 -1862 451146 -1626
rect 451382 -1862 510826 -1626
rect 511062 -1862 511146 -1626
rect 511382 -1862 570826 -1626
rect 571062 -1862 571146 -1626
rect 571382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 4546 -2266
rect 4782 -2502 4866 -2266
rect 5102 -2502 64546 -2266
rect 64782 -2502 64866 -2266
rect 65102 -2502 124546 -2266
rect 124782 -2502 124866 -2266
rect 125102 -2502 184546 -2266
rect 184782 -2502 184866 -2266
rect 185102 -2502 244546 -2266
rect 244782 -2502 244866 -2266
rect 245102 -2502 304546 -2266
rect 304782 -2502 304866 -2266
rect 305102 -2502 364546 -2266
rect 364782 -2502 364866 -2266
rect 365102 -2502 424546 -2266
rect 424782 -2502 424866 -2266
rect 425102 -2502 484546 -2266
rect 484782 -2502 484866 -2266
rect 485102 -2502 544546 -2266
rect 544782 -2502 544866 -2266
rect 545102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 4546 -2586
rect 4782 -2822 4866 -2586
rect 5102 -2822 64546 -2586
rect 64782 -2822 64866 -2586
rect 65102 -2822 124546 -2586
rect 124782 -2822 124866 -2586
rect 125102 -2822 184546 -2586
rect 184782 -2822 184866 -2586
rect 185102 -2822 244546 -2586
rect 244782 -2822 244866 -2586
rect 245102 -2822 304546 -2586
rect 304782 -2822 304866 -2586
rect 305102 -2822 364546 -2586
rect 364782 -2822 364866 -2586
rect 365102 -2822 424546 -2586
rect 424782 -2822 424866 -2586
rect 425102 -2822 484546 -2586
rect 484782 -2822 484866 -2586
rect 485102 -2822 544546 -2586
rect 544782 -2822 544866 -2586
rect 545102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 34546 -3226
rect 34782 -3462 34866 -3226
rect 35102 -3462 94546 -3226
rect 94782 -3462 94866 -3226
rect 95102 -3462 154546 -3226
rect 154782 -3462 154866 -3226
rect 155102 -3462 214546 -3226
rect 214782 -3462 214866 -3226
rect 215102 -3462 274546 -3226
rect 274782 -3462 274866 -3226
rect 275102 -3462 334546 -3226
rect 334782 -3462 334866 -3226
rect 335102 -3462 394546 -3226
rect 394782 -3462 394866 -3226
rect 395102 -3462 454546 -3226
rect 454782 -3462 454866 -3226
rect 455102 -3462 514546 -3226
rect 514782 -3462 514866 -3226
rect 515102 -3462 574546 -3226
rect 574782 -3462 574866 -3226
rect 575102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 34546 -3546
rect 34782 -3782 34866 -3546
rect 35102 -3782 94546 -3546
rect 94782 -3782 94866 -3546
rect 95102 -3782 154546 -3546
rect 154782 -3782 154866 -3546
rect 155102 -3782 214546 -3546
rect 214782 -3782 214866 -3546
rect 215102 -3782 274546 -3546
rect 274782 -3782 274866 -3546
rect 275102 -3782 334546 -3546
rect 334782 -3782 334866 -3546
rect 335102 -3782 394546 -3546
rect 394782 -3782 394866 -3546
rect 395102 -3782 454546 -3546
rect 454782 -3782 454866 -3546
rect 455102 -3782 514546 -3546
rect 514782 -3782 514866 -3546
rect 515102 -3782 574546 -3546
rect 574782 -3782 574866 -3546
rect 575102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 8266 -4186
rect 8502 -4422 8586 -4186
rect 8822 -4422 68266 -4186
rect 68502 -4422 68586 -4186
rect 68822 -4422 128266 -4186
rect 128502 -4422 128586 -4186
rect 128822 -4422 188266 -4186
rect 188502 -4422 188586 -4186
rect 188822 -4422 248266 -4186
rect 248502 -4422 248586 -4186
rect 248822 -4422 308266 -4186
rect 308502 -4422 308586 -4186
rect 308822 -4422 368266 -4186
rect 368502 -4422 368586 -4186
rect 368822 -4422 428266 -4186
rect 428502 -4422 428586 -4186
rect 428822 -4422 488266 -4186
rect 488502 -4422 488586 -4186
rect 488822 -4422 548266 -4186
rect 548502 -4422 548586 -4186
rect 548822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 8266 -4506
rect 8502 -4742 8586 -4506
rect 8822 -4742 68266 -4506
rect 68502 -4742 68586 -4506
rect 68822 -4742 128266 -4506
rect 128502 -4742 128586 -4506
rect 128822 -4742 188266 -4506
rect 188502 -4742 188586 -4506
rect 188822 -4742 248266 -4506
rect 248502 -4742 248586 -4506
rect 248822 -4742 308266 -4506
rect 308502 -4742 308586 -4506
rect 308822 -4742 368266 -4506
rect 368502 -4742 368586 -4506
rect 368822 -4742 428266 -4506
rect 428502 -4742 428586 -4506
rect 428822 -4742 488266 -4506
rect 488502 -4742 488586 -4506
rect 488822 -4742 548266 -4506
rect 548502 -4742 548586 -4506
rect 548822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 38266 -5146
rect 38502 -5382 38586 -5146
rect 38822 -5382 98266 -5146
rect 98502 -5382 98586 -5146
rect 98822 -5382 158266 -5146
rect 158502 -5382 158586 -5146
rect 158822 -5382 218266 -5146
rect 218502 -5382 218586 -5146
rect 218822 -5382 278266 -5146
rect 278502 -5382 278586 -5146
rect 278822 -5382 338266 -5146
rect 338502 -5382 338586 -5146
rect 338822 -5382 398266 -5146
rect 398502 -5382 398586 -5146
rect 398822 -5382 458266 -5146
rect 458502 -5382 458586 -5146
rect 458822 -5382 518266 -5146
rect 518502 -5382 518586 -5146
rect 518822 -5382 578266 -5146
rect 578502 -5382 578586 -5146
rect 578822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 38266 -5466
rect 38502 -5702 38586 -5466
rect 38822 -5702 98266 -5466
rect 98502 -5702 98586 -5466
rect 98822 -5702 158266 -5466
rect 158502 -5702 158586 -5466
rect 158822 -5702 218266 -5466
rect 218502 -5702 218586 -5466
rect 218822 -5702 278266 -5466
rect 278502 -5702 278586 -5466
rect 278822 -5702 338266 -5466
rect 338502 -5702 338586 -5466
rect 338822 -5702 398266 -5466
rect 398502 -5702 398586 -5466
rect 398822 -5702 458266 -5466
rect 458502 -5702 458586 -5466
rect 458822 -5702 518266 -5466
rect 518502 -5702 518586 -5466
rect 518822 -5702 578266 -5466
rect 578502 -5702 578586 -5466
rect 578822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 11986 -6106
rect 12222 -6342 12306 -6106
rect 12542 -6342 71986 -6106
rect 72222 -6342 72306 -6106
rect 72542 -6342 131986 -6106
rect 132222 -6342 132306 -6106
rect 132542 -6342 191986 -6106
rect 192222 -6342 192306 -6106
rect 192542 -6342 251986 -6106
rect 252222 -6342 252306 -6106
rect 252542 -6342 311986 -6106
rect 312222 -6342 312306 -6106
rect 312542 -6342 371986 -6106
rect 372222 -6342 372306 -6106
rect 372542 -6342 431986 -6106
rect 432222 -6342 432306 -6106
rect 432542 -6342 491986 -6106
rect 492222 -6342 492306 -6106
rect 492542 -6342 551986 -6106
rect 552222 -6342 552306 -6106
rect 552542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 11986 -6426
rect 12222 -6662 12306 -6426
rect 12542 -6662 71986 -6426
rect 72222 -6662 72306 -6426
rect 72542 -6662 131986 -6426
rect 132222 -6662 132306 -6426
rect 132542 -6662 191986 -6426
rect 192222 -6662 192306 -6426
rect 192542 -6662 251986 -6426
rect 252222 -6662 252306 -6426
rect 252542 -6662 311986 -6426
rect 312222 -6662 312306 -6426
rect 312542 -6662 371986 -6426
rect 372222 -6662 372306 -6426
rect 372542 -6662 431986 -6426
rect 432222 -6662 432306 -6426
rect 432542 -6662 491986 -6426
rect 492222 -6662 492306 -6426
rect 492542 -6662 551986 -6426
rect 552222 -6662 552306 -6426
rect 552542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 41986 -7066
rect 42222 -7302 42306 -7066
rect 42542 -7302 101986 -7066
rect 102222 -7302 102306 -7066
rect 102542 -7302 161986 -7066
rect 162222 -7302 162306 -7066
rect 162542 -7302 221986 -7066
rect 222222 -7302 222306 -7066
rect 222542 -7302 281986 -7066
rect 282222 -7302 282306 -7066
rect 282542 -7302 341986 -7066
rect 342222 -7302 342306 -7066
rect 342542 -7302 401986 -7066
rect 402222 -7302 402306 -7066
rect 402542 -7302 461986 -7066
rect 462222 -7302 462306 -7066
rect 462542 -7302 521986 -7066
rect 522222 -7302 522306 -7066
rect 522542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 41986 -7386
rect 42222 -7622 42306 -7386
rect 42542 -7622 101986 -7386
rect 102222 -7622 102306 -7386
rect 102542 -7622 161986 -7386
rect 162222 -7622 162306 -7386
rect 162542 -7622 221986 -7386
rect 222222 -7622 222306 -7386
rect 222542 -7622 281986 -7386
rect 282222 -7622 282306 -7386
rect 282542 -7622 341986 -7386
rect 342222 -7622 342306 -7386
rect 342542 -7622 401986 -7386
rect 402222 -7622 402306 -7386
rect 402542 -7622 461986 -7386
rect 462222 -7622 462306 -7386
rect 462542 -7622 521986 -7386
rect 522222 -7622 522306 -7386
rect 522542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use to_ALU_opt_TMR_KP_Voter  TMR_ALU
timestamp 1641133681
transform 1 0 200000 0 1 200000
box 0 0 50151 52295
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 1866 586890 2486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 61866 586890 62486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 121866 586890 122486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 181866 586890 182486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 241866 586890 242486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 301866 586890 302486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 361866 586890 362486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 421866 586890 422486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 481866 586890 482486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 541866 586890 542486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 601866 586890 602486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 661866 586890 662486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 240794 -1894 241414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 794 -1894 1414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 60794 -1894 61414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 120794 -1894 121414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 180794 -1894 181414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 240794 254295 241414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 300794 -1894 301414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 360794 -1894 361414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 420794 -1894 421414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 480794 -1894 481414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 540794 -1894 541414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 5586 588810 6206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 65586 588810 66206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 125586 588810 126206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 185586 588810 186206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 245586 588810 246206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 305586 588810 306206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 365586 588810 366206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 425586 588810 426206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 485586 588810 486206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 545586 588810 546206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 605586 588810 606206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 665586 588810 666206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 244514 -3814 245134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 4514 -3814 5134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 64514 -3814 65134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 124514 -3814 125134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 184514 -3814 185134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 244514 254295 245134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 304514 -3814 305134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 364514 -3814 365134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 424514 -3814 425134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 484514 -3814 485134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 544514 -3814 545134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 9306 590730 9926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 69306 590730 69926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 129306 590730 129926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 189306 590730 189926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 249306 590730 249926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 309306 590730 309926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 369306 590730 369926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 429306 590730 429926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 489306 590730 489926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 549306 590730 549926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 609306 590730 609926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 669306 590730 669926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 248234 -5734 248854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 8234 -5734 8854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 68234 -5734 68854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 128234 -5734 128854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 188234 -5734 188854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 248234 254295 248854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 308234 -5734 308854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 368234 -5734 368854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 428234 -5734 428854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 488234 -5734 488854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 548234 -5734 548854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 13026 592650 13646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 73026 592650 73646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 133026 592650 133646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 193026 592650 193646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 253026 592650 253646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 313026 592650 313646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 373026 592650 373646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 433026 592650 433646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 493026 592650 493646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 553026 592650 553646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 613026 592650 613646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 673026 592650 673646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 251954 -7654 252574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 11954 -7654 12574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 71954 -7654 72574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 131954 -7654 132574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 191954 -7654 192574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 251954 254295 252574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 311954 -7654 312574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 371954 -7654 372574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 431954 -7654 432574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 491954 -7654 492574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 551954 -7654 552574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 39306 590730 39926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 99306 590730 99926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 159306 590730 159926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 219306 590730 219926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 279306 590730 279926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 339306 590730 339926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 399306 590730 399926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 459306 590730 459926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 519306 590730 519926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 579306 590730 579926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 639306 590730 639926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 699306 590730 699926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 218234 -5734 218854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 38234 -5734 38854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 98234 -5734 98854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 158234 -5734 158854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 218234 254295 218854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 278234 -5734 278854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 338234 -5734 338854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 398234 -5734 398854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 458234 -5734 458854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 518234 -5734 518854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 578234 -5734 578854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 43026 592650 43646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 103026 592650 103646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 163026 592650 163646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 223026 592650 223646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 283026 592650 283646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 343026 592650 343646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 403026 592650 403646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 463026 592650 463646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 523026 592650 523646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 583026 592650 583646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 643026 592650 643646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 221954 -7654 222574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 41954 -7654 42574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 101954 -7654 102574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 161954 -7654 162574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 221954 254295 222574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 281954 -7654 282574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 341954 -7654 342574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 401954 -7654 402574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 461954 -7654 462574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 521954 -7654 522574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 31866 586890 32486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 91866 586890 92486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 151866 586890 152486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 211866 586890 212486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 271866 586890 272486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 331866 586890 332486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 391866 586890 392486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 451866 586890 452486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 511866 586890 512486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 571866 586890 572486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 631866 586890 632486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 691866 586890 692486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 210794 -1894 211414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 30794 -1894 31414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 90794 -1894 91414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 150794 -1894 151414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 210794 254295 211414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 270794 -1894 271414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 330794 -1894 331414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 390794 -1894 391414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 450794 -1894 451414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 510794 -1894 511414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 570794 -1894 571414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 35586 588810 36206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 95586 588810 96206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 155586 588810 156206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 215586 588810 216206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 275586 588810 276206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 335586 588810 336206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 395586 588810 396206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 455586 588810 456206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 515586 588810 516206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 575586 588810 576206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 635586 588810 636206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 695586 588810 696206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 214514 -3814 215134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 34514 -3814 35134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 94514 -3814 95134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 154514 -3814 155134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 214514 254295 215134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 274514 -3814 275134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 334514 -3814 335134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 394514 -3814 395134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 454514 -3814 455134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 514514 -3814 515134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 574514 -3814 575134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
